assign W_R_STAGE_LUT[0] = 16'd256;
assign W_I_STAGE_LUT[0] = 16'd0;
assign W_R_STAGE_LUT[1] = 16'd256;
assign W_I_STAGE_LUT[1] = -16'd6;
assign W_R_STAGE_LUT[2] = 16'd256;
assign W_I_STAGE_LUT[2] = -16'd13;
assign W_R_STAGE_LUT[3] = 16'd255;
assign W_I_STAGE_LUT[3] = -16'd19;
assign W_R_STAGE_LUT[4] = 16'd255;
assign W_I_STAGE_LUT[4] = -16'd25;
assign W_R_STAGE_LUT[5] = 16'd254;
assign W_I_STAGE_LUT[5] = -16'd31;
assign W_R_STAGE_LUT[6] = 16'd253;
assign W_I_STAGE_LUT[6] = -16'd38;
assign W_R_STAGE_LUT[7] = 16'd252;
assign W_I_STAGE_LUT[7] = -16'd44;
assign W_R_STAGE_LUT[8] = 16'd251;
assign W_I_STAGE_LUT[8] = -16'd50;
assign W_R_STAGE_LUT[9] = 16'd250;
assign W_I_STAGE_LUT[9] = -16'd56;
assign W_R_STAGE_LUT[10] = 16'd248;
assign W_I_STAGE_LUT[10] = -16'd62;
assign W_R_STAGE_LUT[11] = 16'd247;
assign W_I_STAGE_LUT[11] = -16'd68;
assign W_R_STAGE_LUT[12] = 16'd245;
assign W_I_STAGE_LUT[12] = -16'd74;
assign W_R_STAGE_LUT[13] = 16'd243;
assign W_I_STAGE_LUT[13] = -16'd80;
assign W_R_STAGE_LUT[14] = 16'd241;
assign W_I_STAGE_LUT[14] = -16'd86;
assign W_R_STAGE_LUT[15] = 16'd239;
assign W_I_STAGE_LUT[15] = -16'd92;
assign W_R_STAGE_LUT[16] = 16'd237;
assign W_I_STAGE_LUT[16] = -16'd98;
assign W_R_STAGE_LUT[17] = 16'd234;
assign W_I_STAGE_LUT[17] = -16'd104;
assign W_R_STAGE_LUT[18] = 16'd231;
assign W_I_STAGE_LUT[18] = -16'd109;
assign W_R_STAGE_LUT[19] = 16'd229;
assign W_I_STAGE_LUT[19] = -16'd115;
assign W_R_STAGE_LUT[20] = 16'd226;
assign W_I_STAGE_LUT[20] = -16'd121;
assign W_R_STAGE_LUT[21] = 16'd223;
assign W_I_STAGE_LUT[21] = -16'd126;
assign W_R_STAGE_LUT[22] = 16'd220;
assign W_I_STAGE_LUT[22] = -16'd132;
assign W_R_STAGE_LUT[23] = 16'd216;
assign W_I_STAGE_LUT[23] = -16'd137;
assign W_R_STAGE_LUT[24] = 16'd213;
assign W_I_STAGE_LUT[24] = -16'd142;
assign W_R_STAGE_LUT[25] = 16'd209;
assign W_I_STAGE_LUT[25] = -16'd147;
assign W_R_STAGE_LUT[26] = 16'd206;
assign W_I_STAGE_LUT[26] = -16'd152;
assign W_R_STAGE_LUT[27] = 16'd202;
assign W_I_STAGE_LUT[27] = -16'd157;
assign W_R_STAGE_LUT[28] = 16'd198;
assign W_I_STAGE_LUT[28] = -16'd162;
assign W_R_STAGE_LUT[29] = 16'd194;
assign W_I_STAGE_LUT[29] = -16'd167;
assign W_R_STAGE_LUT[30] = 16'd190;
assign W_I_STAGE_LUT[30] = -16'd172;
assign W_R_STAGE_LUT[31] = 16'd185;
assign W_I_STAGE_LUT[31] = -16'd177;
assign W_R_STAGE_LUT[32] = 16'd181;
assign W_I_STAGE_LUT[32] = -16'd181;
assign W_R_STAGE_LUT[33] = 16'd177;
assign W_I_STAGE_LUT[33] = -16'd185;
assign W_R_STAGE_LUT[34] = 16'd172;
assign W_I_STAGE_LUT[34] = -16'd190;
assign W_R_STAGE_LUT[35] = 16'd167;
assign W_I_STAGE_LUT[35] = -16'd194;
assign W_R_STAGE_LUT[36] = 16'd162;
assign W_I_STAGE_LUT[36] = -16'd198;
assign W_R_STAGE_LUT[37] = 16'd157;
assign W_I_STAGE_LUT[37] = -16'd202;
assign W_R_STAGE_LUT[38] = 16'd152;
assign W_I_STAGE_LUT[38] = -16'd206;
assign W_R_STAGE_LUT[39] = 16'd147;
assign W_I_STAGE_LUT[39] = -16'd209;
assign W_R_STAGE_LUT[40] = 16'd142;
assign W_I_STAGE_LUT[40] = -16'd213;
assign W_R_STAGE_LUT[41] = 16'd137;
assign W_I_STAGE_LUT[41] = -16'd216;
assign W_R_STAGE_LUT[42] = 16'd132;
assign W_I_STAGE_LUT[42] = -16'd220;
assign W_R_STAGE_LUT[43] = 16'd126;
assign W_I_STAGE_LUT[43] = -16'd223;
assign W_R_STAGE_LUT[44] = 16'd121;
assign W_I_STAGE_LUT[44] = -16'd226;
assign W_R_STAGE_LUT[45] = 16'd115;
assign W_I_STAGE_LUT[45] = -16'd229;
assign W_R_STAGE_LUT[46] = 16'd109;
assign W_I_STAGE_LUT[46] = -16'd231;
assign W_R_STAGE_LUT[47] = 16'd104;
assign W_I_STAGE_LUT[47] = -16'd234;
assign W_R_STAGE_LUT[48] = 16'd98;
assign W_I_STAGE_LUT[48] = -16'd237;
assign W_R_STAGE_LUT[49] = 16'd92;
assign W_I_STAGE_LUT[49] = -16'd239;
assign W_R_STAGE_LUT[50] = 16'd86;
assign W_I_STAGE_LUT[50] = -16'd241;
assign W_R_STAGE_LUT[51] = 16'd80;
assign W_I_STAGE_LUT[51] = -16'd243;
assign W_R_STAGE_LUT[52] = 16'd74;
assign W_I_STAGE_LUT[52] = -16'd245;
assign W_R_STAGE_LUT[53] = 16'd68;
assign W_I_STAGE_LUT[53] = -16'd247;
assign W_R_STAGE_LUT[54] = 16'd62;
assign W_I_STAGE_LUT[54] = -16'd248;
assign W_R_STAGE_LUT[55] = 16'd56;
assign W_I_STAGE_LUT[55] = -16'd250;
assign W_R_STAGE_LUT[56] = 16'd50;
assign W_I_STAGE_LUT[56] = -16'd251;
assign W_R_STAGE_LUT[57] = 16'd44;
assign W_I_STAGE_LUT[57] = -16'd252;
assign W_R_STAGE_LUT[58] = 16'd38;
assign W_I_STAGE_LUT[58] = -16'd253;
assign W_R_STAGE_LUT[59] = 16'd31;
assign W_I_STAGE_LUT[59] = -16'd254;
assign W_R_STAGE_LUT[60] = 16'd25;
assign W_I_STAGE_LUT[60] = -16'd255;
assign W_R_STAGE_LUT[61] = 16'd19;
assign W_I_STAGE_LUT[61] = -16'd255;
assign W_R_STAGE_LUT[62] = 16'd13;
assign W_I_STAGE_LUT[62] = -16'd256;
assign W_R_STAGE_LUT[63] = 16'd6;
assign W_I_STAGE_LUT[63] = -16'd256;
assign W_R_STAGE_LUT[64] = 16'd0;
assign W_I_STAGE_LUT[64] = -16'd256;
assign W_R_STAGE_LUT[65] = -16'd6;
assign W_I_STAGE_LUT[65] = -16'd256;
assign W_R_STAGE_LUT[66] = -16'd13;
assign W_I_STAGE_LUT[66] = -16'd256;
assign W_R_STAGE_LUT[67] = -16'd19;
assign W_I_STAGE_LUT[67] = -16'd255;
assign W_R_STAGE_LUT[68] = -16'd25;
assign W_I_STAGE_LUT[68] = -16'd255;
assign W_R_STAGE_LUT[69] = -16'd31;
assign W_I_STAGE_LUT[69] = -16'd254;
assign W_R_STAGE_LUT[70] = -16'd38;
assign W_I_STAGE_LUT[70] = -16'd253;
assign W_R_STAGE_LUT[71] = -16'd44;
assign W_I_STAGE_LUT[71] = -16'd252;
assign W_R_STAGE_LUT[72] = -16'd50;
assign W_I_STAGE_LUT[72] = -16'd251;
assign W_R_STAGE_LUT[73] = -16'd56;
assign W_I_STAGE_LUT[73] = -16'd250;
assign W_R_STAGE_LUT[74] = -16'd62;
assign W_I_STAGE_LUT[74] = -16'd248;
assign W_R_STAGE_LUT[75] = -16'd68;
assign W_I_STAGE_LUT[75] = -16'd247;
assign W_R_STAGE_LUT[76] = -16'd74;
assign W_I_STAGE_LUT[76] = -16'd245;
assign W_R_STAGE_LUT[77] = -16'd80;
assign W_I_STAGE_LUT[77] = -16'd243;
assign W_R_STAGE_LUT[78] = -16'd86;
assign W_I_STAGE_LUT[78] = -16'd241;
assign W_R_STAGE_LUT[79] = -16'd92;
assign W_I_STAGE_LUT[79] = -16'd239;
assign W_R_STAGE_LUT[80] = -16'd98;
assign W_I_STAGE_LUT[80] = -16'd237;
assign W_R_STAGE_LUT[81] = -16'd104;
assign W_I_STAGE_LUT[81] = -16'd234;
assign W_R_STAGE_LUT[82] = -16'd109;
assign W_I_STAGE_LUT[82] = -16'd231;
assign W_R_STAGE_LUT[83] = -16'd115;
assign W_I_STAGE_LUT[83] = -16'd229;
assign W_R_STAGE_LUT[84] = -16'd121;
assign W_I_STAGE_LUT[84] = -16'd226;
assign W_R_STAGE_LUT[85] = -16'd126;
assign W_I_STAGE_LUT[85] = -16'd223;
assign W_R_STAGE_LUT[86] = -16'd132;
assign W_I_STAGE_LUT[86] = -16'd220;
assign W_R_STAGE_LUT[87] = -16'd137;
assign W_I_STAGE_LUT[87] = -16'd216;
assign W_R_STAGE_LUT[88] = -16'd142;
assign W_I_STAGE_LUT[88] = -16'd213;
assign W_R_STAGE_LUT[89] = -16'd147;
assign W_I_STAGE_LUT[89] = -16'd209;
assign W_R_STAGE_LUT[90] = -16'd152;
assign W_I_STAGE_LUT[90] = -16'd206;
assign W_R_STAGE_LUT[91] = -16'd157;
assign W_I_STAGE_LUT[91] = -16'd202;
assign W_R_STAGE_LUT[92] = -16'd162;
assign W_I_STAGE_LUT[92] = -16'd198;
assign W_R_STAGE_LUT[93] = -16'd167;
assign W_I_STAGE_LUT[93] = -16'd194;
assign W_R_STAGE_LUT[94] = -16'd172;
assign W_I_STAGE_LUT[94] = -16'd190;
assign W_R_STAGE_LUT[95] = -16'd177;
assign W_I_STAGE_LUT[95] = -16'd185;
assign W_R_STAGE_LUT[96] = -16'd181;
assign W_I_STAGE_LUT[96] = -16'd181;
assign W_R_STAGE_LUT[97] = -16'd185;
assign W_I_STAGE_LUT[97] = -16'd177;
assign W_R_STAGE_LUT[98] = -16'd190;
assign W_I_STAGE_LUT[98] = -16'd172;
assign W_R_STAGE_LUT[99] = -16'd194;
assign W_I_STAGE_LUT[99] = -16'd167;
assign W_R_STAGE_LUT[100] = -16'd198;
assign W_I_STAGE_LUT[100] = -16'd162;
assign W_R_STAGE_LUT[101] = -16'd202;
assign W_I_STAGE_LUT[101] = -16'd157;
assign W_R_STAGE_LUT[102] = -16'd206;
assign W_I_STAGE_LUT[102] = -16'd152;
assign W_R_STAGE_LUT[103] = -16'd209;
assign W_I_STAGE_LUT[103] = -16'd147;
assign W_R_STAGE_LUT[104] = -16'd213;
assign W_I_STAGE_LUT[104] = -16'd142;
assign W_R_STAGE_LUT[105] = -16'd216;
assign W_I_STAGE_LUT[105] = -16'd137;
assign W_R_STAGE_LUT[106] = -16'd220;
assign W_I_STAGE_LUT[106] = -16'd132;
assign W_R_STAGE_LUT[107] = -16'd223;
assign W_I_STAGE_LUT[107] = -16'd126;
assign W_R_STAGE_LUT[108] = -16'd226;
assign W_I_STAGE_LUT[108] = -16'd121;
assign W_R_STAGE_LUT[109] = -16'd229;
assign W_I_STAGE_LUT[109] = -16'd115;
assign W_R_STAGE_LUT[110] = -16'd231;
assign W_I_STAGE_LUT[110] = -16'd109;
assign W_R_STAGE_LUT[111] = -16'd234;
assign W_I_STAGE_LUT[111] = -16'd104;
assign W_R_STAGE_LUT[112] = -16'd237;
assign W_I_STAGE_LUT[112] = -16'd98;
assign W_R_STAGE_LUT[113] = -16'd239;
assign W_I_STAGE_LUT[113] = -16'd92;
assign W_R_STAGE_LUT[114] = -16'd241;
assign W_I_STAGE_LUT[114] = -16'd86;
assign W_R_STAGE_LUT[115] = -16'd243;
assign W_I_STAGE_LUT[115] = -16'd80;
assign W_R_STAGE_LUT[116] = -16'd245;
assign W_I_STAGE_LUT[116] = -16'd74;
assign W_R_STAGE_LUT[117] = -16'd247;
assign W_I_STAGE_LUT[117] = -16'd68;
assign W_R_STAGE_LUT[118] = -16'd248;
assign W_I_STAGE_LUT[118] = -16'd62;
assign W_R_STAGE_LUT[119] = -16'd250;
assign W_I_STAGE_LUT[119] = -16'd56;
assign W_R_STAGE_LUT[120] = -16'd251;
assign W_I_STAGE_LUT[120] = -16'd50;
assign W_R_STAGE_LUT[121] = -16'd252;
assign W_I_STAGE_LUT[121] = -16'd44;
assign W_R_STAGE_LUT[122] = -16'd253;
assign W_I_STAGE_LUT[122] = -16'd38;
assign W_R_STAGE_LUT[123] = -16'd254;
assign W_I_STAGE_LUT[123] = -16'd31;
assign W_R_STAGE_LUT[124] = -16'd255;
assign W_I_STAGE_LUT[124] = -16'd25;
assign W_R_STAGE_LUT[125] = -16'd255;
assign W_I_STAGE_LUT[125] = -16'd19;
assign W_R_STAGE_LUT[126] = -16'd256;
assign W_I_STAGE_LUT[126] = -16'd13;
assign W_R_STAGE_LUT[127] = -16'd256;
assign W_I_STAGE_LUT[127] = -16'd6;
