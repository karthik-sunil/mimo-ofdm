assign W_R_STAGE_LUT[0] = 16'd256;
assign W_I_STAGE_LUT[0] = 16'd0;
assign W_R_STAGE_LUT[1] = 16'd256;
assign W_I_STAGE_LUT[1] = 16'd0;
assign W_R_STAGE_LUT[2] = 16'd256;
assign W_I_STAGE_LUT[2] = -16'd1;
assign W_R_STAGE_LUT[3] = 16'd256;
assign W_I_STAGE_LUT[3] = -16'd1;
assign W_R_STAGE_LUT[4] = 16'd256;
assign W_I_STAGE_LUT[4] = -16'd2;
assign W_R_STAGE_LUT[5] = 16'd256;
assign W_I_STAGE_LUT[5] = -16'd2;
assign W_R_STAGE_LUT[6] = 16'd256;
assign W_I_STAGE_LUT[6] = -16'd2;
assign W_R_STAGE_LUT[7] = 16'd256;
assign W_I_STAGE_LUT[7] = -16'd3;
assign W_R_STAGE_LUT[8] = 16'd256;
assign W_I_STAGE_LUT[8] = -16'd3;
assign W_R_STAGE_LUT[9] = 16'd256;
assign W_I_STAGE_LUT[9] = -16'd4;
assign W_R_STAGE_LUT[10] = 16'd256;
assign W_I_STAGE_LUT[10] = -16'd4;
assign W_R_STAGE_LUT[11] = 16'd256;
assign W_I_STAGE_LUT[11] = -16'd4;
assign W_R_STAGE_LUT[12] = 16'd256;
assign W_I_STAGE_LUT[12] = -16'd5;
assign W_R_STAGE_LUT[13] = 16'd256;
assign W_I_STAGE_LUT[13] = -16'd5;
assign W_R_STAGE_LUT[14] = 16'd256;
assign W_I_STAGE_LUT[14] = -16'd5;
assign W_R_STAGE_LUT[15] = 16'd256;
assign W_I_STAGE_LUT[15] = -16'd6;
assign W_R_STAGE_LUT[16] = 16'd256;
assign W_I_STAGE_LUT[16] = -16'd6;
assign W_R_STAGE_LUT[17] = 16'd256;
assign W_I_STAGE_LUT[17] = -16'd7;
assign W_R_STAGE_LUT[18] = 16'd256;
assign W_I_STAGE_LUT[18] = -16'd7;
assign W_R_STAGE_LUT[19] = 16'd256;
assign W_I_STAGE_LUT[19] = -16'd7;
assign W_R_STAGE_LUT[20] = 16'd256;
assign W_I_STAGE_LUT[20] = -16'd8;
assign W_R_STAGE_LUT[21] = 16'd256;
assign W_I_STAGE_LUT[21] = -16'd8;
assign W_R_STAGE_LUT[22] = 16'd256;
assign W_I_STAGE_LUT[22] = -16'd9;
assign W_R_STAGE_LUT[23] = 16'd256;
assign W_I_STAGE_LUT[23] = -16'd9;
assign W_R_STAGE_LUT[24] = 16'd256;
assign W_I_STAGE_LUT[24] = -16'd9;
assign W_R_STAGE_LUT[25] = 16'd256;
assign W_I_STAGE_LUT[25] = -16'd10;
assign W_R_STAGE_LUT[26] = 16'd256;
assign W_I_STAGE_LUT[26] = -16'd10;
assign W_R_STAGE_LUT[27] = 16'd256;
assign W_I_STAGE_LUT[27] = -16'd11;
assign W_R_STAGE_LUT[28] = 16'd256;
assign W_I_STAGE_LUT[28] = -16'd11;
assign W_R_STAGE_LUT[29] = 16'd256;
assign W_I_STAGE_LUT[29] = -16'd11;
assign W_R_STAGE_LUT[30] = 16'd256;
assign W_I_STAGE_LUT[30] = -16'd12;
assign W_R_STAGE_LUT[31] = 16'd256;
assign W_I_STAGE_LUT[31] = -16'd12;
assign W_R_STAGE_LUT[32] = 16'd256;
assign W_I_STAGE_LUT[32] = -16'd13;
assign W_R_STAGE_LUT[33] = 16'd256;
assign W_I_STAGE_LUT[33] = -16'd13;
assign W_R_STAGE_LUT[34] = 16'd256;
assign W_I_STAGE_LUT[34] = -16'd13;
assign W_R_STAGE_LUT[35] = 16'd256;
assign W_I_STAGE_LUT[35] = -16'd14;
assign W_R_STAGE_LUT[36] = 16'd256;
assign W_I_STAGE_LUT[36] = -16'd14;
assign W_R_STAGE_LUT[37] = 16'd256;
assign W_I_STAGE_LUT[37] = -16'd15;
assign W_R_STAGE_LUT[38] = 16'd256;
assign W_I_STAGE_LUT[38] = -16'd15;
assign W_R_STAGE_LUT[39] = 16'd256;
assign W_I_STAGE_LUT[39] = -16'd15;
assign W_R_STAGE_LUT[40] = 16'd256;
assign W_I_STAGE_LUT[40] = -16'd16;
assign W_R_STAGE_LUT[41] = 16'd255;
assign W_I_STAGE_LUT[41] = -16'd16;
assign W_R_STAGE_LUT[42] = 16'd255;
assign W_I_STAGE_LUT[42] = -16'd16;
assign W_R_STAGE_LUT[43] = 16'd255;
assign W_I_STAGE_LUT[43] = -16'd17;
assign W_R_STAGE_LUT[44] = 16'd255;
assign W_I_STAGE_LUT[44] = -16'd17;
assign W_R_STAGE_LUT[45] = 16'd255;
assign W_I_STAGE_LUT[45] = -16'd18;
assign W_R_STAGE_LUT[46] = 16'd255;
assign W_I_STAGE_LUT[46] = -16'd18;
assign W_R_STAGE_LUT[47] = 16'd255;
assign W_I_STAGE_LUT[47] = -16'd18;
assign W_R_STAGE_LUT[48] = 16'd255;
assign W_I_STAGE_LUT[48] = -16'd19;
assign W_R_STAGE_LUT[49] = 16'd255;
assign W_I_STAGE_LUT[49] = -16'd19;
assign W_R_STAGE_LUT[50] = 16'd255;
assign W_I_STAGE_LUT[50] = -16'd20;
assign W_R_STAGE_LUT[51] = 16'd255;
assign W_I_STAGE_LUT[51] = -16'd20;
assign W_R_STAGE_LUT[52] = 16'd255;
assign W_I_STAGE_LUT[52] = -16'd20;
assign W_R_STAGE_LUT[53] = 16'd255;
assign W_I_STAGE_LUT[53] = -16'd21;
assign W_R_STAGE_LUT[54] = 16'd255;
assign W_I_STAGE_LUT[54] = -16'd21;
assign W_R_STAGE_LUT[55] = 16'd255;
assign W_I_STAGE_LUT[55] = -16'd22;
assign W_R_STAGE_LUT[56] = 16'd255;
assign W_I_STAGE_LUT[56] = -16'd22;
assign W_R_STAGE_LUT[57] = 16'd255;
assign W_I_STAGE_LUT[57] = -16'd22;
assign W_R_STAGE_LUT[58] = 16'd255;
assign W_I_STAGE_LUT[58] = -16'd23;
assign W_R_STAGE_LUT[59] = 16'd255;
assign W_I_STAGE_LUT[59] = -16'd23;
assign W_R_STAGE_LUT[60] = 16'd255;
assign W_I_STAGE_LUT[60] = -16'd24;
assign W_R_STAGE_LUT[61] = 16'd255;
assign W_I_STAGE_LUT[61] = -16'd24;
assign W_R_STAGE_LUT[62] = 16'd255;
assign W_I_STAGE_LUT[62] = -16'd24;
assign W_R_STAGE_LUT[63] = 16'd255;
assign W_I_STAGE_LUT[63] = -16'd25;
assign W_R_STAGE_LUT[64] = 16'd255;
assign W_I_STAGE_LUT[64] = -16'd25;
assign W_R_STAGE_LUT[65] = 16'd255;
assign W_I_STAGE_LUT[65] = -16'd25;
assign W_R_STAGE_LUT[66] = 16'd255;
assign W_I_STAGE_LUT[66] = -16'd26;
assign W_R_STAGE_LUT[67] = 16'd255;
assign W_I_STAGE_LUT[67] = -16'd26;
assign W_R_STAGE_LUT[68] = 16'd255;
assign W_I_STAGE_LUT[68] = -16'd27;
assign W_R_STAGE_LUT[69] = 16'd255;
assign W_I_STAGE_LUT[69] = -16'd27;
assign W_R_STAGE_LUT[70] = 16'd255;
assign W_I_STAGE_LUT[70] = -16'd27;
assign W_R_STAGE_LUT[71] = 16'd254;
assign W_I_STAGE_LUT[71] = -16'd28;
assign W_R_STAGE_LUT[72] = 16'd254;
assign W_I_STAGE_LUT[72] = -16'd28;
assign W_R_STAGE_LUT[73] = 16'd254;
assign W_I_STAGE_LUT[73] = -16'd29;
assign W_R_STAGE_LUT[74] = 16'd254;
assign W_I_STAGE_LUT[74] = -16'd29;
assign W_R_STAGE_LUT[75] = 16'd254;
assign W_I_STAGE_LUT[75] = -16'd29;
assign W_R_STAGE_LUT[76] = 16'd254;
assign W_I_STAGE_LUT[76] = -16'd30;
assign W_R_STAGE_LUT[77] = 16'd254;
assign W_I_STAGE_LUT[77] = -16'd30;
assign W_R_STAGE_LUT[78] = 16'd254;
assign W_I_STAGE_LUT[78] = -16'd31;
assign W_R_STAGE_LUT[79] = 16'd254;
assign W_I_STAGE_LUT[79] = -16'd31;
assign W_R_STAGE_LUT[80] = 16'd254;
assign W_I_STAGE_LUT[80] = -16'd31;
assign W_R_STAGE_LUT[81] = 16'd254;
assign W_I_STAGE_LUT[81] = -16'd32;
assign W_R_STAGE_LUT[82] = 16'd254;
assign W_I_STAGE_LUT[82] = -16'd32;
assign W_R_STAGE_LUT[83] = 16'd254;
assign W_I_STAGE_LUT[83] = -16'd33;
assign W_R_STAGE_LUT[84] = 16'd254;
assign W_I_STAGE_LUT[84] = -16'd33;
assign W_R_STAGE_LUT[85] = 16'd254;
assign W_I_STAGE_LUT[85] = -16'd33;
assign W_R_STAGE_LUT[86] = 16'd254;
assign W_I_STAGE_LUT[86] = -16'd34;
assign W_R_STAGE_LUT[87] = 16'd254;
assign W_I_STAGE_LUT[87] = -16'd34;
assign W_R_STAGE_LUT[88] = 16'd254;
assign W_I_STAGE_LUT[88] = -16'd34;
assign W_R_STAGE_LUT[89] = 16'd254;
assign W_I_STAGE_LUT[89] = -16'd35;
assign W_R_STAGE_LUT[90] = 16'd254;
assign W_I_STAGE_LUT[90] = -16'd35;
assign W_R_STAGE_LUT[91] = 16'd254;
assign W_I_STAGE_LUT[91] = -16'd36;
assign W_R_STAGE_LUT[92] = 16'd253;
assign W_I_STAGE_LUT[92] = -16'd36;
assign W_R_STAGE_LUT[93] = 16'd253;
assign W_I_STAGE_LUT[93] = -16'd36;
assign W_R_STAGE_LUT[94] = 16'd253;
assign W_I_STAGE_LUT[94] = -16'd37;
assign W_R_STAGE_LUT[95] = 16'd253;
assign W_I_STAGE_LUT[95] = -16'd37;
assign W_R_STAGE_LUT[96] = 16'd253;
assign W_I_STAGE_LUT[96] = -16'd38;
assign W_R_STAGE_LUT[97] = 16'd253;
assign W_I_STAGE_LUT[97] = -16'd38;
assign W_R_STAGE_LUT[98] = 16'd253;
assign W_I_STAGE_LUT[98] = -16'd38;
assign W_R_STAGE_LUT[99] = 16'd253;
assign W_I_STAGE_LUT[99] = -16'd39;
assign W_R_STAGE_LUT[100] = 16'd253;
assign W_I_STAGE_LUT[100] = -16'd39;
assign W_R_STAGE_LUT[101] = 16'd253;
assign W_I_STAGE_LUT[101] = -16'd40;
assign W_R_STAGE_LUT[102] = 16'd253;
assign W_I_STAGE_LUT[102] = -16'd40;
assign W_R_STAGE_LUT[103] = 16'd253;
assign W_I_STAGE_LUT[103] = -16'd40;
assign W_R_STAGE_LUT[104] = 16'd253;
assign W_I_STAGE_LUT[104] = -16'd41;
assign W_R_STAGE_LUT[105] = 16'd253;
assign W_I_STAGE_LUT[105] = -16'd41;
assign W_R_STAGE_LUT[106] = 16'd253;
assign W_I_STAGE_LUT[106] = -16'd41;
assign W_R_STAGE_LUT[107] = 16'd253;
assign W_I_STAGE_LUT[107] = -16'd42;
assign W_R_STAGE_LUT[108] = 16'd252;
assign W_I_STAGE_LUT[108] = -16'd42;
assign W_R_STAGE_LUT[109] = 16'd252;
assign W_I_STAGE_LUT[109] = -16'd43;
assign W_R_STAGE_LUT[110] = 16'd252;
assign W_I_STAGE_LUT[110] = -16'd43;
assign W_R_STAGE_LUT[111] = 16'd252;
assign W_I_STAGE_LUT[111] = -16'd43;
assign W_R_STAGE_LUT[112] = 16'd252;
assign W_I_STAGE_LUT[112] = -16'd44;
assign W_R_STAGE_LUT[113] = 16'd252;
assign W_I_STAGE_LUT[113] = -16'd44;
assign W_R_STAGE_LUT[114] = 16'd252;
assign W_I_STAGE_LUT[114] = -16'd45;
assign W_R_STAGE_LUT[115] = 16'd252;
assign W_I_STAGE_LUT[115] = -16'd45;
assign W_R_STAGE_LUT[116] = 16'd252;
assign W_I_STAGE_LUT[116] = -16'd45;
assign W_R_STAGE_LUT[117] = 16'd252;
assign W_I_STAGE_LUT[117] = -16'd46;
assign W_R_STAGE_LUT[118] = 16'd252;
assign W_I_STAGE_LUT[118] = -16'd46;
assign W_R_STAGE_LUT[119] = 16'd252;
assign W_I_STAGE_LUT[119] = -16'd46;
assign W_R_STAGE_LUT[120] = 16'd252;
assign W_I_STAGE_LUT[120] = -16'd47;
assign W_R_STAGE_LUT[121] = 16'd252;
assign W_I_STAGE_LUT[121] = -16'd47;
assign W_R_STAGE_LUT[122] = 16'd252;
assign W_I_STAGE_LUT[122] = -16'd48;
assign W_R_STAGE_LUT[123] = 16'd251;
assign W_I_STAGE_LUT[123] = -16'd48;
assign W_R_STAGE_LUT[124] = 16'd251;
assign W_I_STAGE_LUT[124] = -16'd48;
assign W_R_STAGE_LUT[125] = 16'd251;
assign W_I_STAGE_LUT[125] = -16'd49;
assign W_R_STAGE_LUT[126] = 16'd251;
assign W_I_STAGE_LUT[126] = -16'd49;
assign W_R_STAGE_LUT[127] = 16'd251;
assign W_I_STAGE_LUT[127] = -16'd50;
assign W_R_STAGE_LUT[128] = 16'd251;
assign W_I_STAGE_LUT[128] = -16'd50;
assign W_R_STAGE_LUT[129] = 16'd251;
assign W_I_STAGE_LUT[129] = -16'd50;
assign W_R_STAGE_LUT[130] = 16'd251;
assign W_I_STAGE_LUT[130] = -16'd51;
assign W_R_STAGE_LUT[131] = 16'd251;
assign W_I_STAGE_LUT[131] = -16'd51;
assign W_R_STAGE_LUT[132] = 16'd251;
assign W_I_STAGE_LUT[132] = -16'd51;
assign W_R_STAGE_LUT[133] = 16'd251;
assign W_I_STAGE_LUT[133] = -16'd52;
assign W_R_STAGE_LUT[134] = 16'd251;
assign W_I_STAGE_LUT[134] = -16'd52;
assign W_R_STAGE_LUT[135] = 16'd251;
assign W_I_STAGE_LUT[135] = -16'd53;
assign W_R_STAGE_LUT[136] = 16'd250;
assign W_I_STAGE_LUT[136] = -16'd53;
assign W_R_STAGE_LUT[137] = 16'd250;
assign W_I_STAGE_LUT[137] = -16'd53;
assign W_R_STAGE_LUT[138] = 16'd250;
assign W_I_STAGE_LUT[138] = -16'd54;
assign W_R_STAGE_LUT[139] = 16'd250;
assign W_I_STAGE_LUT[139] = -16'd54;
assign W_R_STAGE_LUT[140] = 16'd250;
assign W_I_STAGE_LUT[140] = -16'd55;
assign W_R_STAGE_LUT[141] = 16'd250;
assign W_I_STAGE_LUT[141] = -16'd55;
assign W_R_STAGE_LUT[142] = 16'd250;
assign W_I_STAGE_LUT[142] = -16'd55;
assign W_R_STAGE_LUT[143] = 16'd250;
assign W_I_STAGE_LUT[143] = -16'd56;
assign W_R_STAGE_LUT[144] = 16'd250;
assign W_I_STAGE_LUT[144] = -16'd56;
assign W_R_STAGE_LUT[145] = 16'd250;
assign W_I_STAGE_LUT[145] = -16'd56;
assign W_R_STAGE_LUT[146] = 16'd250;
assign W_I_STAGE_LUT[146] = -16'd57;
assign W_R_STAGE_LUT[147] = 16'd250;
assign W_I_STAGE_LUT[147] = -16'd57;
assign W_R_STAGE_LUT[148] = 16'd249;
assign W_I_STAGE_LUT[148] = -16'd58;
assign W_R_STAGE_LUT[149] = 16'd249;
assign W_I_STAGE_LUT[149] = -16'd58;
assign W_R_STAGE_LUT[150] = 16'd249;
assign W_I_STAGE_LUT[150] = -16'd58;
assign W_R_STAGE_LUT[151] = 16'd249;
assign W_I_STAGE_LUT[151] = -16'd59;
assign W_R_STAGE_LUT[152] = 16'd249;
assign W_I_STAGE_LUT[152] = -16'd59;
assign W_R_STAGE_LUT[153] = 16'd249;
assign W_I_STAGE_LUT[153] = -16'd60;
assign W_R_STAGE_LUT[154] = 16'd249;
assign W_I_STAGE_LUT[154] = -16'd60;
assign W_R_STAGE_LUT[155] = 16'd249;
assign W_I_STAGE_LUT[155] = -16'd60;
assign W_R_STAGE_LUT[156] = 16'd249;
assign W_I_STAGE_LUT[156] = -16'd61;
assign W_R_STAGE_LUT[157] = 16'd249;
assign W_I_STAGE_LUT[157] = -16'd61;
assign W_R_STAGE_LUT[158] = 16'd249;
assign W_I_STAGE_LUT[158] = -16'd61;
assign W_R_STAGE_LUT[159] = 16'd248;
assign W_I_STAGE_LUT[159] = -16'd62;
assign W_R_STAGE_LUT[160] = 16'd248;
assign W_I_STAGE_LUT[160] = -16'd62;
assign W_R_STAGE_LUT[161] = 16'd248;
assign W_I_STAGE_LUT[161] = -16'd63;
assign W_R_STAGE_LUT[162] = 16'd248;
assign W_I_STAGE_LUT[162] = -16'd63;
assign W_R_STAGE_LUT[163] = 16'd248;
assign W_I_STAGE_LUT[163] = -16'd63;
assign W_R_STAGE_LUT[164] = 16'd248;
assign W_I_STAGE_LUT[164] = -16'd64;
assign W_R_STAGE_LUT[165] = 16'd248;
assign W_I_STAGE_LUT[165] = -16'd64;
assign W_R_STAGE_LUT[166] = 16'd248;
assign W_I_STAGE_LUT[166] = -16'd64;
assign W_R_STAGE_LUT[167] = 16'd248;
assign W_I_STAGE_LUT[167] = -16'd65;
assign W_R_STAGE_LUT[168] = 16'd248;
assign W_I_STAGE_LUT[168] = -16'd65;
assign W_R_STAGE_LUT[169] = 16'd247;
assign W_I_STAGE_LUT[169] = -16'd66;
assign W_R_STAGE_LUT[170] = 16'd247;
assign W_I_STAGE_LUT[170] = -16'd66;
assign W_R_STAGE_LUT[171] = 16'd247;
assign W_I_STAGE_LUT[171] = -16'd66;
assign W_R_STAGE_LUT[172] = 16'd247;
assign W_I_STAGE_LUT[172] = -16'd67;
assign W_R_STAGE_LUT[173] = 16'd247;
assign W_I_STAGE_LUT[173] = -16'd67;
assign W_R_STAGE_LUT[174] = 16'd247;
assign W_I_STAGE_LUT[174] = -16'd68;
assign W_R_STAGE_LUT[175] = 16'd247;
assign W_I_STAGE_LUT[175] = -16'd68;
assign W_R_STAGE_LUT[176] = 16'd247;
assign W_I_STAGE_LUT[176] = -16'd68;
assign W_R_STAGE_LUT[177] = 16'd247;
assign W_I_STAGE_LUT[177] = -16'd69;
assign W_R_STAGE_LUT[178] = 16'd247;
assign W_I_STAGE_LUT[178] = -16'd69;
assign W_R_STAGE_LUT[179] = 16'd246;
assign W_I_STAGE_LUT[179] = -16'd69;
assign W_R_STAGE_LUT[180] = 16'd246;
assign W_I_STAGE_LUT[180] = -16'd70;
assign W_R_STAGE_LUT[181] = 16'd246;
assign W_I_STAGE_LUT[181] = -16'd70;
assign W_R_STAGE_LUT[182] = 16'd246;
assign W_I_STAGE_LUT[182] = -16'd71;
assign W_R_STAGE_LUT[183] = 16'd246;
assign W_I_STAGE_LUT[183] = -16'd71;
assign W_R_STAGE_LUT[184] = 16'd246;
assign W_I_STAGE_LUT[184] = -16'd71;
assign W_R_STAGE_LUT[185] = 16'd246;
assign W_I_STAGE_LUT[185] = -16'd72;
assign W_R_STAGE_LUT[186] = 16'd246;
assign W_I_STAGE_LUT[186] = -16'd72;
assign W_R_STAGE_LUT[187] = 16'd246;
assign W_I_STAGE_LUT[187] = -16'd72;
assign W_R_STAGE_LUT[188] = 16'd245;
assign W_I_STAGE_LUT[188] = -16'd73;
assign W_R_STAGE_LUT[189] = 16'd245;
assign W_I_STAGE_LUT[189] = -16'd73;
assign W_R_STAGE_LUT[190] = 16'd245;
assign W_I_STAGE_LUT[190] = -16'd74;
assign W_R_STAGE_LUT[191] = 16'd245;
assign W_I_STAGE_LUT[191] = -16'd74;
assign W_R_STAGE_LUT[192] = 16'd245;
assign W_I_STAGE_LUT[192] = -16'd74;
assign W_R_STAGE_LUT[193] = 16'd245;
assign W_I_STAGE_LUT[193] = -16'd75;
assign W_R_STAGE_LUT[194] = 16'd245;
assign W_I_STAGE_LUT[194] = -16'd75;
assign W_R_STAGE_LUT[195] = 16'd245;
assign W_I_STAGE_LUT[195] = -16'd75;
assign W_R_STAGE_LUT[196] = 16'd245;
assign W_I_STAGE_LUT[196] = -16'd76;
assign W_R_STAGE_LUT[197] = 16'd244;
assign W_I_STAGE_LUT[197] = -16'd76;
assign W_R_STAGE_LUT[198] = 16'd244;
assign W_I_STAGE_LUT[198] = -16'd77;
assign W_R_STAGE_LUT[199] = 16'd244;
assign W_I_STAGE_LUT[199] = -16'd77;
assign W_R_STAGE_LUT[200] = 16'd244;
assign W_I_STAGE_LUT[200] = -16'd77;
assign W_R_STAGE_LUT[201] = 16'd244;
assign W_I_STAGE_LUT[201] = -16'd78;
assign W_R_STAGE_LUT[202] = 16'd244;
assign W_I_STAGE_LUT[202] = -16'd78;
assign W_R_STAGE_LUT[203] = 16'd244;
assign W_I_STAGE_LUT[203] = -16'd78;
assign W_R_STAGE_LUT[204] = 16'd244;
assign W_I_STAGE_LUT[204] = -16'd79;
assign W_R_STAGE_LUT[205] = 16'd243;
assign W_I_STAGE_LUT[205] = -16'd79;
assign W_R_STAGE_LUT[206] = 16'd243;
assign W_I_STAGE_LUT[206] = -16'd80;
assign W_R_STAGE_LUT[207] = 16'd243;
assign W_I_STAGE_LUT[207] = -16'd80;
assign W_R_STAGE_LUT[208] = 16'd243;
assign W_I_STAGE_LUT[208] = -16'd80;
assign W_R_STAGE_LUT[209] = 16'd243;
assign W_I_STAGE_LUT[209] = -16'd81;
assign W_R_STAGE_LUT[210] = 16'd243;
assign W_I_STAGE_LUT[210] = -16'd81;
assign W_R_STAGE_LUT[211] = 16'd243;
assign W_I_STAGE_LUT[211] = -16'd81;
assign W_R_STAGE_LUT[212] = 16'd243;
assign W_I_STAGE_LUT[212] = -16'd82;
assign W_R_STAGE_LUT[213] = 16'd242;
assign W_I_STAGE_LUT[213] = -16'd82;
assign W_R_STAGE_LUT[214] = 16'd242;
assign W_I_STAGE_LUT[214] = -16'd83;
assign W_R_STAGE_LUT[215] = 16'd242;
assign W_I_STAGE_LUT[215] = -16'd83;
assign W_R_STAGE_LUT[216] = 16'd242;
assign W_I_STAGE_LUT[216] = -16'd83;
assign W_R_STAGE_LUT[217] = 16'd242;
assign W_I_STAGE_LUT[217] = -16'd84;
assign W_R_STAGE_LUT[218] = 16'd242;
assign W_I_STAGE_LUT[218] = -16'd84;
assign W_R_STAGE_LUT[219] = 16'd242;
assign W_I_STAGE_LUT[219] = -16'd84;
assign W_R_STAGE_LUT[220] = 16'd242;
assign W_I_STAGE_LUT[220] = -16'd85;
assign W_R_STAGE_LUT[221] = 16'd241;
assign W_I_STAGE_LUT[221] = -16'd85;
assign W_R_STAGE_LUT[222] = 16'd241;
assign W_I_STAGE_LUT[222] = -16'd86;
assign W_R_STAGE_LUT[223] = 16'd241;
assign W_I_STAGE_LUT[223] = -16'd86;
assign W_R_STAGE_LUT[224] = 16'd241;
assign W_I_STAGE_LUT[224] = -16'd86;
assign W_R_STAGE_LUT[225] = 16'd241;
assign W_I_STAGE_LUT[225] = -16'd87;
assign W_R_STAGE_LUT[226] = 16'd241;
assign W_I_STAGE_LUT[226] = -16'd87;
assign W_R_STAGE_LUT[227] = 16'd241;
assign W_I_STAGE_LUT[227] = -16'd87;
assign W_R_STAGE_LUT[228] = 16'd241;
assign W_I_STAGE_LUT[228] = -16'd88;
assign W_R_STAGE_LUT[229] = 16'd240;
assign W_I_STAGE_LUT[229] = -16'd88;
assign W_R_STAGE_LUT[230] = 16'd240;
assign W_I_STAGE_LUT[230] = -16'd88;
assign W_R_STAGE_LUT[231] = 16'd240;
assign W_I_STAGE_LUT[231] = -16'd89;
assign W_R_STAGE_LUT[232] = 16'd240;
assign W_I_STAGE_LUT[232] = -16'd89;
assign W_R_STAGE_LUT[233] = 16'd240;
assign W_I_STAGE_LUT[233] = -16'd90;
assign W_R_STAGE_LUT[234] = 16'd240;
assign W_I_STAGE_LUT[234] = -16'd90;
assign W_R_STAGE_LUT[235] = 16'd240;
assign W_I_STAGE_LUT[235] = -16'd90;
assign W_R_STAGE_LUT[236] = 16'd239;
assign W_I_STAGE_LUT[236] = -16'd91;
assign W_R_STAGE_LUT[237] = 16'd239;
assign W_I_STAGE_LUT[237] = -16'd91;
assign W_R_STAGE_LUT[238] = 16'd239;
assign W_I_STAGE_LUT[238] = -16'd91;
assign W_R_STAGE_LUT[239] = 16'd239;
assign W_I_STAGE_LUT[239] = -16'd92;
assign W_R_STAGE_LUT[240] = 16'd239;
assign W_I_STAGE_LUT[240] = -16'd92;
assign W_R_STAGE_LUT[241] = 16'd239;
assign W_I_STAGE_LUT[241] = -16'd92;
assign W_R_STAGE_LUT[242] = 16'd239;
assign W_I_STAGE_LUT[242] = -16'd93;
assign W_R_STAGE_LUT[243] = 16'd238;
assign W_I_STAGE_LUT[243] = -16'd93;
assign W_R_STAGE_LUT[244] = 16'd238;
assign W_I_STAGE_LUT[244] = -16'd94;
assign W_R_STAGE_LUT[245] = 16'd238;
assign W_I_STAGE_LUT[245] = -16'd94;
assign W_R_STAGE_LUT[246] = 16'd238;
assign W_I_STAGE_LUT[246] = -16'd94;
assign W_R_STAGE_LUT[247] = 16'd238;
assign W_I_STAGE_LUT[247] = -16'd95;
assign W_R_STAGE_LUT[248] = 16'd238;
assign W_I_STAGE_LUT[248] = -16'd95;
assign W_R_STAGE_LUT[249] = 16'd238;
assign W_I_STAGE_LUT[249] = -16'd95;
assign W_R_STAGE_LUT[250] = 16'd237;
assign W_I_STAGE_LUT[250] = -16'd96;
assign W_R_STAGE_LUT[251] = 16'd237;
assign W_I_STAGE_LUT[251] = -16'd96;
assign W_R_STAGE_LUT[252] = 16'd237;
assign W_I_STAGE_LUT[252] = -16'd97;
assign W_R_STAGE_LUT[253] = 16'd237;
assign W_I_STAGE_LUT[253] = -16'd97;
assign W_R_STAGE_LUT[254] = 16'd237;
assign W_I_STAGE_LUT[254] = -16'd97;
assign W_R_STAGE_LUT[255] = 16'd237;
assign W_I_STAGE_LUT[255] = -16'd98;
assign W_R_STAGE_LUT[256] = 16'd237;
assign W_I_STAGE_LUT[256] = -16'd98;
assign W_R_STAGE_LUT[257] = 16'd236;
assign W_I_STAGE_LUT[257] = -16'd98;
assign W_R_STAGE_LUT[258] = 16'd236;
assign W_I_STAGE_LUT[258] = -16'd99;
assign W_R_STAGE_LUT[259] = 16'd236;
assign W_I_STAGE_LUT[259] = -16'd99;
assign W_R_STAGE_LUT[260] = 16'd236;
assign W_I_STAGE_LUT[260] = -16'd99;
assign W_R_STAGE_LUT[261] = 16'd236;
assign W_I_STAGE_LUT[261] = -16'd100;
assign W_R_STAGE_LUT[262] = 16'd236;
assign W_I_STAGE_LUT[262] = -16'd100;
assign W_R_STAGE_LUT[263] = 16'd235;
assign W_I_STAGE_LUT[263] = -16'd101;
assign W_R_STAGE_LUT[264] = 16'd235;
assign W_I_STAGE_LUT[264] = -16'd101;
assign W_R_STAGE_LUT[265] = 16'd235;
assign W_I_STAGE_LUT[265] = -16'd101;
assign W_R_STAGE_LUT[266] = 16'd235;
assign W_I_STAGE_LUT[266] = -16'd102;
assign W_R_STAGE_LUT[267] = 16'd235;
assign W_I_STAGE_LUT[267] = -16'd102;
assign W_R_STAGE_LUT[268] = 16'd235;
assign W_I_STAGE_LUT[268] = -16'd102;
assign W_R_STAGE_LUT[269] = 16'd235;
assign W_I_STAGE_LUT[269] = -16'd103;
assign W_R_STAGE_LUT[270] = 16'd234;
assign W_I_STAGE_LUT[270] = -16'd103;
assign W_R_STAGE_LUT[271] = 16'd234;
assign W_I_STAGE_LUT[271] = -16'd103;
assign W_R_STAGE_LUT[272] = 16'd234;
assign W_I_STAGE_LUT[272] = -16'd104;
assign W_R_STAGE_LUT[273] = 16'd234;
assign W_I_STAGE_LUT[273] = -16'd104;
assign W_R_STAGE_LUT[274] = 16'd234;
assign W_I_STAGE_LUT[274] = -16'd104;
assign W_R_STAGE_LUT[275] = 16'd234;
assign W_I_STAGE_LUT[275] = -16'd105;
assign W_R_STAGE_LUT[276] = 16'd233;
assign W_I_STAGE_LUT[276] = -16'd105;
assign W_R_STAGE_LUT[277] = 16'd233;
assign W_I_STAGE_LUT[277] = -16'd106;
assign W_R_STAGE_LUT[278] = 16'd233;
assign W_I_STAGE_LUT[278] = -16'd106;
assign W_R_STAGE_LUT[279] = 16'd233;
assign W_I_STAGE_LUT[279] = -16'd106;
assign W_R_STAGE_LUT[280] = 16'd233;
assign W_I_STAGE_LUT[280] = -16'd107;
assign W_R_STAGE_LUT[281] = 16'd233;
assign W_I_STAGE_LUT[281] = -16'd107;
assign W_R_STAGE_LUT[282] = 16'd232;
assign W_I_STAGE_LUT[282] = -16'd107;
assign W_R_STAGE_LUT[283] = 16'd232;
assign W_I_STAGE_LUT[283] = -16'd108;
assign W_R_STAGE_LUT[284] = 16'd232;
assign W_I_STAGE_LUT[284] = -16'd108;
assign W_R_STAGE_LUT[285] = 16'd232;
assign W_I_STAGE_LUT[285] = -16'd108;
assign W_R_STAGE_LUT[286] = 16'd232;
assign W_I_STAGE_LUT[286] = -16'd109;
assign W_R_STAGE_LUT[287] = 16'd232;
assign W_I_STAGE_LUT[287] = -16'd109;
assign W_R_STAGE_LUT[288] = 16'd231;
assign W_I_STAGE_LUT[288] = -16'd109;
assign W_R_STAGE_LUT[289] = 16'd231;
assign W_I_STAGE_LUT[289] = -16'd110;
assign W_R_STAGE_LUT[290] = 16'd231;
assign W_I_STAGE_LUT[290] = -16'd110;
assign W_R_STAGE_LUT[291] = 16'd231;
assign W_I_STAGE_LUT[291] = -16'd111;
assign W_R_STAGE_LUT[292] = 16'd231;
assign W_I_STAGE_LUT[292] = -16'd111;
assign W_R_STAGE_LUT[293] = 16'd231;
assign W_I_STAGE_LUT[293] = -16'd111;
assign W_R_STAGE_LUT[294] = 16'd230;
assign W_I_STAGE_LUT[294] = -16'd112;
assign W_R_STAGE_LUT[295] = 16'd230;
assign W_I_STAGE_LUT[295] = -16'd112;
assign W_R_STAGE_LUT[296] = 16'd230;
assign W_I_STAGE_LUT[296] = -16'd112;
assign W_R_STAGE_LUT[297] = 16'd230;
assign W_I_STAGE_LUT[297] = -16'd113;
assign W_R_STAGE_LUT[298] = 16'd230;
assign W_I_STAGE_LUT[298] = -16'd113;
assign W_R_STAGE_LUT[299] = 16'd230;
assign W_I_STAGE_LUT[299] = -16'd113;
assign W_R_STAGE_LUT[300] = 16'd229;
assign W_I_STAGE_LUT[300] = -16'd114;
assign W_R_STAGE_LUT[301] = 16'd229;
assign W_I_STAGE_LUT[301] = -16'd114;
assign W_R_STAGE_LUT[302] = 16'd229;
assign W_I_STAGE_LUT[302] = -16'd114;
assign W_R_STAGE_LUT[303] = 16'd229;
assign W_I_STAGE_LUT[303] = -16'd115;
assign W_R_STAGE_LUT[304] = 16'd229;
assign W_I_STAGE_LUT[304] = -16'd115;
assign W_R_STAGE_LUT[305] = 16'd228;
assign W_I_STAGE_LUT[305] = -16'd115;
assign W_R_STAGE_LUT[306] = 16'd228;
assign W_I_STAGE_LUT[306] = -16'd116;
assign W_R_STAGE_LUT[307] = 16'd228;
assign W_I_STAGE_LUT[307] = -16'd116;
assign W_R_STAGE_LUT[308] = 16'd228;
assign W_I_STAGE_LUT[308] = -16'd117;
assign W_R_STAGE_LUT[309] = 16'd228;
assign W_I_STAGE_LUT[309] = -16'd117;
assign W_R_STAGE_LUT[310] = 16'd228;
assign W_I_STAGE_LUT[310] = -16'd117;
assign W_R_STAGE_LUT[311] = 16'd227;
assign W_I_STAGE_LUT[311] = -16'd118;
assign W_R_STAGE_LUT[312] = 16'd227;
assign W_I_STAGE_LUT[312] = -16'd118;
assign W_R_STAGE_LUT[313] = 16'd227;
assign W_I_STAGE_LUT[313] = -16'd118;
assign W_R_STAGE_LUT[314] = 16'd227;
assign W_I_STAGE_LUT[314] = -16'd119;
assign W_R_STAGE_LUT[315] = 16'd227;
assign W_I_STAGE_LUT[315] = -16'd119;
assign W_R_STAGE_LUT[316] = 16'd227;
assign W_I_STAGE_LUT[316] = -16'd119;
assign W_R_STAGE_LUT[317] = 16'd226;
assign W_I_STAGE_LUT[317] = -16'd120;
assign W_R_STAGE_LUT[318] = 16'd226;
assign W_I_STAGE_LUT[318] = -16'd120;
assign W_R_STAGE_LUT[319] = 16'd226;
assign W_I_STAGE_LUT[319] = -16'd120;
assign W_R_STAGE_LUT[320] = 16'd226;
assign W_I_STAGE_LUT[320] = -16'd121;
assign W_R_STAGE_LUT[321] = 16'd226;
assign W_I_STAGE_LUT[321] = -16'd121;
assign W_R_STAGE_LUT[322] = 16'd225;
assign W_I_STAGE_LUT[322] = -16'd121;
assign W_R_STAGE_LUT[323] = 16'd225;
assign W_I_STAGE_LUT[323] = -16'd122;
assign W_R_STAGE_LUT[324] = 16'd225;
assign W_I_STAGE_LUT[324] = -16'd122;
assign W_R_STAGE_LUT[325] = 16'd225;
assign W_I_STAGE_LUT[325] = -16'd122;
assign W_R_STAGE_LUT[326] = 16'd225;
assign W_I_STAGE_LUT[326] = -16'd123;
assign W_R_STAGE_LUT[327] = 16'd224;
assign W_I_STAGE_LUT[327] = -16'd123;
assign W_R_STAGE_LUT[328] = 16'd224;
assign W_I_STAGE_LUT[328] = -16'd123;
assign W_R_STAGE_LUT[329] = 16'd224;
assign W_I_STAGE_LUT[329] = -16'd124;
assign W_R_STAGE_LUT[330] = 16'd224;
assign W_I_STAGE_LUT[330] = -16'd124;
assign W_R_STAGE_LUT[331] = 16'd224;
assign W_I_STAGE_LUT[331] = -16'd124;
assign W_R_STAGE_LUT[332] = 16'd224;
assign W_I_STAGE_LUT[332] = -16'd125;
assign W_R_STAGE_LUT[333] = 16'd223;
assign W_I_STAGE_LUT[333] = -16'd125;
assign W_R_STAGE_LUT[334] = 16'd223;
assign W_I_STAGE_LUT[334] = -16'd125;
assign W_R_STAGE_LUT[335] = 16'd223;
assign W_I_STAGE_LUT[335] = -16'd126;
assign W_R_STAGE_LUT[336] = 16'd223;
assign W_I_STAGE_LUT[336] = -16'd126;
assign W_R_STAGE_LUT[337] = 16'd223;
assign W_I_STAGE_LUT[337] = -16'd127;
assign W_R_STAGE_LUT[338] = 16'd222;
assign W_I_STAGE_LUT[338] = -16'd127;
assign W_R_STAGE_LUT[339] = 16'd222;
assign W_I_STAGE_LUT[339] = -16'd127;
assign W_R_STAGE_LUT[340] = 16'd222;
assign W_I_STAGE_LUT[340] = -16'd128;
assign W_R_STAGE_LUT[341] = 16'd222;
assign W_I_STAGE_LUT[341] = -16'd128;
assign W_R_STAGE_LUT[342] = 16'd222;
assign W_I_STAGE_LUT[342] = -16'd128;
assign W_R_STAGE_LUT[343] = 16'd221;
assign W_I_STAGE_LUT[343] = -16'd129;
assign W_R_STAGE_LUT[344] = 16'd221;
assign W_I_STAGE_LUT[344] = -16'd129;
assign W_R_STAGE_LUT[345] = 16'd221;
assign W_I_STAGE_LUT[345] = -16'd129;
assign W_R_STAGE_LUT[346] = 16'd221;
assign W_I_STAGE_LUT[346] = -16'd130;
assign W_R_STAGE_LUT[347] = 16'd221;
assign W_I_STAGE_LUT[347] = -16'd130;
assign W_R_STAGE_LUT[348] = 16'd220;
assign W_I_STAGE_LUT[348] = -16'd130;
assign W_R_STAGE_LUT[349] = 16'd220;
assign W_I_STAGE_LUT[349] = -16'd131;
assign W_R_STAGE_LUT[350] = 16'd220;
assign W_I_STAGE_LUT[350] = -16'd131;
assign W_R_STAGE_LUT[351] = 16'd220;
assign W_I_STAGE_LUT[351] = -16'd131;
assign W_R_STAGE_LUT[352] = 16'd220;
assign W_I_STAGE_LUT[352] = -16'd132;
assign W_R_STAGE_LUT[353] = 16'd219;
assign W_I_STAGE_LUT[353] = -16'd132;
assign W_R_STAGE_LUT[354] = 16'd219;
assign W_I_STAGE_LUT[354] = -16'd132;
assign W_R_STAGE_LUT[355] = 16'd219;
assign W_I_STAGE_LUT[355] = -16'd133;
assign W_R_STAGE_LUT[356] = 16'd219;
assign W_I_STAGE_LUT[356] = -16'd133;
assign W_R_STAGE_LUT[357] = 16'd219;
assign W_I_STAGE_LUT[357] = -16'd133;
assign W_R_STAGE_LUT[358] = 16'd218;
assign W_I_STAGE_LUT[358] = -16'd134;
assign W_R_STAGE_LUT[359] = 16'd218;
assign W_I_STAGE_LUT[359] = -16'd134;
assign W_R_STAGE_LUT[360] = 16'd218;
assign W_I_STAGE_LUT[360] = -16'd134;
assign W_R_STAGE_LUT[361] = 16'd218;
assign W_I_STAGE_LUT[361] = -16'd135;
assign W_R_STAGE_LUT[362] = 16'd218;
assign W_I_STAGE_LUT[362] = -16'd135;
assign W_R_STAGE_LUT[363] = 16'd217;
assign W_I_STAGE_LUT[363] = -16'd135;
assign W_R_STAGE_LUT[364] = 16'd217;
assign W_I_STAGE_LUT[364] = -16'd136;
assign W_R_STAGE_LUT[365] = 16'd217;
assign W_I_STAGE_LUT[365] = -16'd136;
assign W_R_STAGE_LUT[366] = 16'd217;
assign W_I_STAGE_LUT[366] = -16'd136;
assign W_R_STAGE_LUT[367] = 16'd216;
assign W_I_STAGE_LUT[367] = -16'd137;
assign W_R_STAGE_LUT[368] = 16'd216;
assign W_I_STAGE_LUT[368] = -16'd137;
assign W_R_STAGE_LUT[369] = 16'd216;
assign W_I_STAGE_LUT[369] = -16'd137;
assign W_R_STAGE_LUT[370] = 16'd216;
assign W_I_STAGE_LUT[370] = -16'd138;
assign W_R_STAGE_LUT[371] = 16'd216;
assign W_I_STAGE_LUT[371] = -16'd138;
assign W_R_STAGE_LUT[372] = 16'd215;
assign W_I_STAGE_LUT[372] = -16'd138;
assign W_R_STAGE_LUT[373] = 16'd215;
assign W_I_STAGE_LUT[373] = -16'd139;
assign W_R_STAGE_LUT[374] = 16'd215;
assign W_I_STAGE_LUT[374] = -16'd139;
assign W_R_STAGE_LUT[375] = 16'd215;
assign W_I_STAGE_LUT[375] = -16'd139;
assign W_R_STAGE_LUT[376] = 16'd215;
assign W_I_STAGE_LUT[376] = -16'd140;
assign W_R_STAGE_LUT[377] = 16'd214;
assign W_I_STAGE_LUT[377] = -16'd140;
assign W_R_STAGE_LUT[378] = 16'd214;
assign W_I_STAGE_LUT[378] = -16'd140;
assign W_R_STAGE_LUT[379] = 16'd214;
assign W_I_STAGE_LUT[379] = -16'd141;
assign W_R_STAGE_LUT[380] = 16'd214;
assign W_I_STAGE_LUT[380] = -16'd141;
assign W_R_STAGE_LUT[381] = 16'd214;
assign W_I_STAGE_LUT[381] = -16'd141;
assign W_R_STAGE_LUT[382] = 16'd213;
assign W_I_STAGE_LUT[382] = -16'd142;
assign W_R_STAGE_LUT[383] = 16'd213;
assign W_I_STAGE_LUT[383] = -16'd142;
assign W_R_STAGE_LUT[384] = 16'd213;
assign W_I_STAGE_LUT[384] = -16'd142;
assign W_R_STAGE_LUT[385] = 16'd213;
assign W_I_STAGE_LUT[385] = -16'd143;
assign W_R_STAGE_LUT[386] = 16'd212;
assign W_I_STAGE_LUT[386] = -16'd143;
assign W_R_STAGE_LUT[387] = 16'd212;
assign W_I_STAGE_LUT[387] = -16'd143;
assign W_R_STAGE_LUT[388] = 16'd212;
assign W_I_STAGE_LUT[388] = -16'd144;
assign W_R_STAGE_LUT[389] = 16'd212;
assign W_I_STAGE_LUT[389] = -16'd144;
assign W_R_STAGE_LUT[390] = 16'd212;
assign W_I_STAGE_LUT[390] = -16'd144;
assign W_R_STAGE_LUT[391] = 16'd211;
assign W_I_STAGE_LUT[391] = -16'd145;
assign W_R_STAGE_LUT[392] = 16'd211;
assign W_I_STAGE_LUT[392] = -16'd145;
assign W_R_STAGE_LUT[393] = 16'd211;
assign W_I_STAGE_LUT[393] = -16'd145;
assign W_R_STAGE_LUT[394] = 16'd211;
assign W_I_STAGE_LUT[394] = -16'd145;
assign W_R_STAGE_LUT[395] = 16'd210;
assign W_I_STAGE_LUT[395] = -16'd146;
assign W_R_STAGE_LUT[396] = 16'd210;
assign W_I_STAGE_LUT[396] = -16'd146;
assign W_R_STAGE_LUT[397] = 16'd210;
assign W_I_STAGE_LUT[397] = -16'd146;
assign W_R_STAGE_LUT[398] = 16'd210;
assign W_I_STAGE_LUT[398] = -16'd147;
assign W_R_STAGE_LUT[399] = 16'd210;
assign W_I_STAGE_LUT[399] = -16'd147;
assign W_R_STAGE_LUT[400] = 16'd209;
assign W_I_STAGE_LUT[400] = -16'd147;
assign W_R_STAGE_LUT[401] = 16'd209;
assign W_I_STAGE_LUT[401] = -16'd148;
assign W_R_STAGE_LUT[402] = 16'd209;
assign W_I_STAGE_LUT[402] = -16'd148;
assign W_R_STAGE_LUT[403] = 16'd209;
assign W_I_STAGE_LUT[403] = -16'd148;
assign W_R_STAGE_LUT[404] = 16'd208;
assign W_I_STAGE_LUT[404] = -16'd149;
assign W_R_STAGE_LUT[405] = 16'd208;
assign W_I_STAGE_LUT[405] = -16'd149;
assign W_R_STAGE_LUT[406] = 16'd208;
assign W_I_STAGE_LUT[406] = -16'd149;
assign W_R_STAGE_LUT[407] = 16'd208;
assign W_I_STAGE_LUT[407] = -16'd150;
assign W_R_STAGE_LUT[408] = 16'd207;
assign W_I_STAGE_LUT[408] = -16'd150;
assign W_R_STAGE_LUT[409] = 16'd207;
assign W_I_STAGE_LUT[409] = -16'd150;
assign W_R_STAGE_LUT[410] = 16'd207;
assign W_I_STAGE_LUT[410] = -16'd151;
assign W_R_STAGE_LUT[411] = 16'd207;
assign W_I_STAGE_LUT[411] = -16'd151;
assign W_R_STAGE_LUT[412] = 16'd207;
assign W_I_STAGE_LUT[412] = -16'd151;
assign W_R_STAGE_LUT[413] = 16'd206;
assign W_I_STAGE_LUT[413] = -16'd152;
assign W_R_STAGE_LUT[414] = 16'd206;
assign W_I_STAGE_LUT[414] = -16'd152;
assign W_R_STAGE_LUT[415] = 16'd206;
assign W_I_STAGE_LUT[415] = -16'd152;
assign W_R_STAGE_LUT[416] = 16'd206;
assign W_I_STAGE_LUT[416] = -16'd152;
assign W_R_STAGE_LUT[417] = 16'd205;
assign W_I_STAGE_LUT[417] = -16'd153;
assign W_R_STAGE_LUT[418] = 16'd205;
assign W_I_STAGE_LUT[418] = -16'd153;
assign W_R_STAGE_LUT[419] = 16'd205;
assign W_I_STAGE_LUT[419] = -16'd153;
assign W_R_STAGE_LUT[420] = 16'd205;
assign W_I_STAGE_LUT[420] = -16'd154;
assign W_R_STAGE_LUT[421] = 16'd204;
assign W_I_STAGE_LUT[421] = -16'd154;
assign W_R_STAGE_LUT[422] = 16'd204;
assign W_I_STAGE_LUT[422] = -16'd154;
assign W_R_STAGE_LUT[423] = 16'd204;
assign W_I_STAGE_LUT[423] = -16'd155;
assign W_R_STAGE_LUT[424] = 16'd204;
assign W_I_STAGE_LUT[424] = -16'd155;
assign W_R_STAGE_LUT[425] = 16'd203;
assign W_I_STAGE_LUT[425] = -16'd155;
assign W_R_STAGE_LUT[426] = 16'd203;
assign W_I_STAGE_LUT[426] = -16'd156;
assign W_R_STAGE_LUT[427] = 16'd203;
assign W_I_STAGE_LUT[427] = -16'd156;
assign W_R_STAGE_LUT[428] = 16'd203;
assign W_I_STAGE_LUT[428] = -16'd156;
assign W_R_STAGE_LUT[429] = 16'd203;
assign W_I_STAGE_LUT[429] = -16'd157;
assign W_R_STAGE_LUT[430] = 16'd202;
assign W_I_STAGE_LUT[430] = -16'd157;
assign W_R_STAGE_LUT[431] = 16'd202;
assign W_I_STAGE_LUT[431] = -16'd157;
assign W_R_STAGE_LUT[432] = 16'd202;
assign W_I_STAGE_LUT[432] = -16'd157;
assign W_R_STAGE_LUT[433] = 16'd202;
assign W_I_STAGE_LUT[433] = -16'd158;
assign W_R_STAGE_LUT[434] = 16'd201;
assign W_I_STAGE_LUT[434] = -16'd158;
assign W_R_STAGE_LUT[435] = 16'd201;
assign W_I_STAGE_LUT[435] = -16'd158;
assign W_R_STAGE_LUT[436] = 16'd201;
assign W_I_STAGE_LUT[436] = -16'd159;
assign W_R_STAGE_LUT[437] = 16'd201;
assign W_I_STAGE_LUT[437] = -16'd159;
assign W_R_STAGE_LUT[438] = 16'd200;
assign W_I_STAGE_LUT[438] = -16'd159;
assign W_R_STAGE_LUT[439] = 16'd200;
assign W_I_STAGE_LUT[439] = -16'd160;
assign W_R_STAGE_LUT[440] = 16'd200;
assign W_I_STAGE_LUT[440] = -16'd160;
assign W_R_STAGE_LUT[441] = 16'd200;
assign W_I_STAGE_LUT[441] = -16'd160;
assign W_R_STAGE_LUT[442] = 16'd199;
assign W_I_STAGE_LUT[442] = -16'd161;
assign W_R_STAGE_LUT[443] = 16'd199;
assign W_I_STAGE_LUT[443] = -16'd161;
assign W_R_STAGE_LUT[444] = 16'd199;
assign W_I_STAGE_LUT[444] = -16'd161;
assign W_R_STAGE_LUT[445] = 16'd199;
assign W_I_STAGE_LUT[445] = -16'd161;
assign W_R_STAGE_LUT[446] = 16'd198;
assign W_I_STAGE_LUT[446] = -16'd162;
assign W_R_STAGE_LUT[447] = 16'd198;
assign W_I_STAGE_LUT[447] = -16'd162;
assign W_R_STAGE_LUT[448] = 16'd198;
assign W_I_STAGE_LUT[448] = -16'd162;
assign W_R_STAGE_LUT[449] = 16'd198;
assign W_I_STAGE_LUT[449] = -16'd163;
assign W_R_STAGE_LUT[450] = 16'd197;
assign W_I_STAGE_LUT[450] = -16'd163;
assign W_R_STAGE_LUT[451] = 16'd197;
assign W_I_STAGE_LUT[451] = -16'd163;
assign W_R_STAGE_LUT[452] = 16'd197;
assign W_I_STAGE_LUT[452] = -16'd164;
assign W_R_STAGE_LUT[453] = 16'd197;
assign W_I_STAGE_LUT[453] = -16'd164;
assign W_R_STAGE_LUT[454] = 16'd196;
assign W_I_STAGE_LUT[454] = -16'd164;
assign W_R_STAGE_LUT[455] = 16'd196;
assign W_I_STAGE_LUT[455] = -16'd165;
assign W_R_STAGE_LUT[456] = 16'd196;
assign W_I_STAGE_LUT[456] = -16'd165;
assign W_R_STAGE_LUT[457] = 16'd196;
assign W_I_STAGE_LUT[457] = -16'd165;
assign W_R_STAGE_LUT[458] = 16'd195;
assign W_I_STAGE_LUT[458] = -16'd165;
assign W_R_STAGE_LUT[459] = 16'd195;
assign W_I_STAGE_LUT[459] = -16'd166;
assign W_R_STAGE_LUT[460] = 16'd195;
assign W_I_STAGE_LUT[460] = -16'd166;
assign W_R_STAGE_LUT[461] = 16'd195;
assign W_I_STAGE_LUT[461] = -16'd166;
assign W_R_STAGE_LUT[462] = 16'd194;
assign W_I_STAGE_LUT[462] = -16'd167;
assign W_R_STAGE_LUT[463] = 16'd194;
assign W_I_STAGE_LUT[463] = -16'd167;
assign W_R_STAGE_LUT[464] = 16'd194;
assign W_I_STAGE_LUT[464] = -16'd167;
assign W_R_STAGE_LUT[465] = 16'd194;
assign W_I_STAGE_LUT[465] = -16'd168;
assign W_R_STAGE_LUT[466] = 16'd193;
assign W_I_STAGE_LUT[466] = -16'd168;
assign W_R_STAGE_LUT[467] = 16'd193;
assign W_I_STAGE_LUT[467] = -16'd168;
assign W_R_STAGE_LUT[468] = 16'd193;
assign W_I_STAGE_LUT[468] = -16'd168;
assign W_R_STAGE_LUT[469] = 16'd193;
assign W_I_STAGE_LUT[469] = -16'd169;
assign W_R_STAGE_LUT[470] = 16'd192;
assign W_I_STAGE_LUT[470] = -16'd169;
assign W_R_STAGE_LUT[471] = 16'd192;
assign W_I_STAGE_LUT[471] = -16'd169;
assign W_R_STAGE_LUT[472] = 16'd192;
assign W_I_STAGE_LUT[472] = -16'd170;
assign W_R_STAGE_LUT[473] = 16'd192;
assign W_I_STAGE_LUT[473] = -16'd170;
assign W_R_STAGE_LUT[474] = 16'd191;
assign W_I_STAGE_LUT[474] = -16'd170;
assign W_R_STAGE_LUT[475] = 16'd191;
assign W_I_STAGE_LUT[475] = -16'd170;
assign W_R_STAGE_LUT[476] = 16'd191;
assign W_I_STAGE_LUT[476] = -16'd171;
assign W_R_STAGE_LUT[477] = 16'd190;
assign W_I_STAGE_LUT[477] = -16'd171;
assign W_R_STAGE_LUT[478] = 16'd190;
assign W_I_STAGE_LUT[478] = -16'd171;
assign W_R_STAGE_LUT[479] = 16'd190;
assign W_I_STAGE_LUT[479] = -16'd172;
assign W_R_STAGE_LUT[480] = 16'd190;
assign W_I_STAGE_LUT[480] = -16'd172;
assign W_R_STAGE_LUT[481] = 16'd189;
assign W_I_STAGE_LUT[481] = -16'd172;
assign W_R_STAGE_LUT[482] = 16'd189;
assign W_I_STAGE_LUT[482] = -16'd173;
assign W_R_STAGE_LUT[483] = 16'd189;
assign W_I_STAGE_LUT[483] = -16'd173;
assign W_R_STAGE_LUT[484] = 16'd189;
assign W_I_STAGE_LUT[484] = -16'd173;
assign W_R_STAGE_LUT[485] = 16'd188;
assign W_I_STAGE_LUT[485] = -16'd173;
assign W_R_STAGE_LUT[486] = 16'd188;
assign W_I_STAGE_LUT[486] = -16'd174;
assign W_R_STAGE_LUT[487] = 16'd188;
assign W_I_STAGE_LUT[487] = -16'd174;
assign W_R_STAGE_LUT[488] = 16'd188;
assign W_I_STAGE_LUT[488] = -16'd174;
assign W_R_STAGE_LUT[489] = 16'd187;
assign W_I_STAGE_LUT[489] = -16'd175;
assign W_R_STAGE_LUT[490] = 16'd187;
assign W_I_STAGE_LUT[490] = -16'd175;
assign W_R_STAGE_LUT[491] = 16'd187;
assign W_I_STAGE_LUT[491] = -16'd175;
assign W_R_STAGE_LUT[492] = 16'd186;
assign W_I_STAGE_LUT[492] = -16'd175;
assign W_R_STAGE_LUT[493] = 16'd186;
assign W_I_STAGE_LUT[493] = -16'd176;
assign W_R_STAGE_LUT[494] = 16'd186;
assign W_I_STAGE_LUT[494] = -16'd176;
assign W_R_STAGE_LUT[495] = 16'd186;
assign W_I_STAGE_LUT[495] = -16'd176;
assign W_R_STAGE_LUT[496] = 16'd185;
assign W_I_STAGE_LUT[496] = -16'd177;
assign W_R_STAGE_LUT[497] = 16'd185;
assign W_I_STAGE_LUT[497] = -16'd177;
assign W_R_STAGE_LUT[498] = 16'd185;
assign W_I_STAGE_LUT[498] = -16'd177;
assign W_R_STAGE_LUT[499] = 16'd185;
assign W_I_STAGE_LUT[499] = -16'd177;
assign W_R_STAGE_LUT[500] = 16'd184;
assign W_I_STAGE_LUT[500] = -16'd178;
assign W_R_STAGE_LUT[501] = 16'd184;
assign W_I_STAGE_LUT[501] = -16'd178;
assign W_R_STAGE_LUT[502] = 16'd184;
assign W_I_STAGE_LUT[502] = -16'd178;
assign W_R_STAGE_LUT[503] = 16'd184;
assign W_I_STAGE_LUT[503] = -16'd179;
assign W_R_STAGE_LUT[504] = 16'd183;
assign W_I_STAGE_LUT[504] = -16'd179;
assign W_R_STAGE_LUT[505] = 16'd183;
assign W_I_STAGE_LUT[505] = -16'd179;
assign W_R_STAGE_LUT[506] = 16'd183;
assign W_I_STAGE_LUT[506] = -16'd179;
assign W_R_STAGE_LUT[507] = 16'd182;
assign W_I_STAGE_LUT[507] = -16'd180;
assign W_R_STAGE_LUT[508] = 16'd182;
assign W_I_STAGE_LUT[508] = -16'd180;
assign W_R_STAGE_LUT[509] = 16'd182;
assign W_I_STAGE_LUT[509] = -16'd180;
assign W_R_STAGE_LUT[510] = 16'd182;
assign W_I_STAGE_LUT[510] = -16'd180;
assign W_R_STAGE_LUT[511] = 16'd181;
assign W_I_STAGE_LUT[511] = -16'd181;
assign W_R_STAGE_LUT[512] = 16'd181;
assign W_I_STAGE_LUT[512] = -16'd181;
assign W_R_STAGE_LUT[513] = 16'd181;
assign W_I_STAGE_LUT[513] = -16'd181;
assign W_R_STAGE_LUT[514] = 16'd180;
assign W_I_STAGE_LUT[514] = -16'd182;
assign W_R_STAGE_LUT[515] = 16'd180;
assign W_I_STAGE_LUT[515] = -16'd182;
assign W_R_STAGE_LUT[516] = 16'd180;
assign W_I_STAGE_LUT[516] = -16'd182;
assign W_R_STAGE_LUT[517] = 16'd180;
assign W_I_STAGE_LUT[517] = -16'd182;
assign W_R_STAGE_LUT[518] = 16'd179;
assign W_I_STAGE_LUT[518] = -16'd183;
assign W_R_STAGE_LUT[519] = 16'd179;
assign W_I_STAGE_LUT[519] = -16'd183;
assign W_R_STAGE_LUT[520] = 16'd179;
assign W_I_STAGE_LUT[520] = -16'd183;
assign W_R_STAGE_LUT[521] = 16'd179;
assign W_I_STAGE_LUT[521] = -16'd184;
assign W_R_STAGE_LUT[522] = 16'd178;
assign W_I_STAGE_LUT[522] = -16'd184;
assign W_R_STAGE_LUT[523] = 16'd178;
assign W_I_STAGE_LUT[523] = -16'd184;
assign W_R_STAGE_LUT[524] = 16'd178;
assign W_I_STAGE_LUT[524] = -16'd184;
assign W_R_STAGE_LUT[525] = 16'd177;
assign W_I_STAGE_LUT[525] = -16'd185;
assign W_R_STAGE_LUT[526] = 16'd177;
assign W_I_STAGE_LUT[526] = -16'd185;
assign W_R_STAGE_LUT[527] = 16'd177;
assign W_I_STAGE_LUT[527] = -16'd185;
assign W_R_STAGE_LUT[528] = 16'd177;
assign W_I_STAGE_LUT[528] = -16'd185;
assign W_R_STAGE_LUT[529] = 16'd176;
assign W_I_STAGE_LUT[529] = -16'd186;
assign W_R_STAGE_LUT[530] = 16'd176;
assign W_I_STAGE_LUT[530] = -16'd186;
assign W_R_STAGE_LUT[531] = 16'd176;
assign W_I_STAGE_LUT[531] = -16'd186;
assign W_R_STAGE_LUT[532] = 16'd175;
assign W_I_STAGE_LUT[532] = -16'd186;
assign W_R_STAGE_LUT[533] = 16'd175;
assign W_I_STAGE_LUT[533] = -16'd187;
assign W_R_STAGE_LUT[534] = 16'd175;
assign W_I_STAGE_LUT[534] = -16'd187;
assign W_R_STAGE_LUT[535] = 16'd175;
assign W_I_STAGE_LUT[535] = -16'd187;
assign W_R_STAGE_LUT[536] = 16'd174;
assign W_I_STAGE_LUT[536] = -16'd188;
assign W_R_STAGE_LUT[537] = 16'd174;
assign W_I_STAGE_LUT[537] = -16'd188;
assign W_R_STAGE_LUT[538] = 16'd174;
assign W_I_STAGE_LUT[538] = -16'd188;
assign W_R_STAGE_LUT[539] = 16'd173;
assign W_I_STAGE_LUT[539] = -16'd188;
assign W_R_STAGE_LUT[540] = 16'd173;
assign W_I_STAGE_LUT[540] = -16'd189;
assign W_R_STAGE_LUT[541] = 16'd173;
assign W_I_STAGE_LUT[541] = -16'd189;
assign W_R_STAGE_LUT[542] = 16'd173;
assign W_I_STAGE_LUT[542] = -16'd189;
assign W_R_STAGE_LUT[543] = 16'd172;
assign W_I_STAGE_LUT[543] = -16'd189;
assign W_R_STAGE_LUT[544] = 16'd172;
assign W_I_STAGE_LUT[544] = -16'd190;
assign W_R_STAGE_LUT[545] = 16'd172;
assign W_I_STAGE_LUT[545] = -16'd190;
assign W_R_STAGE_LUT[546] = 16'd171;
assign W_I_STAGE_LUT[546] = -16'd190;
assign W_R_STAGE_LUT[547] = 16'd171;
assign W_I_STAGE_LUT[547] = -16'd190;
assign W_R_STAGE_LUT[548] = 16'd171;
assign W_I_STAGE_LUT[548] = -16'd191;
assign W_R_STAGE_LUT[549] = 16'd170;
assign W_I_STAGE_LUT[549] = -16'd191;
assign W_R_STAGE_LUT[550] = 16'd170;
assign W_I_STAGE_LUT[550] = -16'd191;
assign W_R_STAGE_LUT[551] = 16'd170;
assign W_I_STAGE_LUT[551] = -16'd192;
assign W_R_STAGE_LUT[552] = 16'd170;
assign W_I_STAGE_LUT[552] = -16'd192;
assign W_R_STAGE_LUT[553] = 16'd169;
assign W_I_STAGE_LUT[553] = -16'd192;
assign W_R_STAGE_LUT[554] = 16'd169;
assign W_I_STAGE_LUT[554] = -16'd192;
assign W_R_STAGE_LUT[555] = 16'd169;
assign W_I_STAGE_LUT[555] = -16'd193;
assign W_R_STAGE_LUT[556] = 16'd168;
assign W_I_STAGE_LUT[556] = -16'd193;
assign W_R_STAGE_LUT[557] = 16'd168;
assign W_I_STAGE_LUT[557] = -16'd193;
assign W_R_STAGE_LUT[558] = 16'd168;
assign W_I_STAGE_LUT[558] = -16'd193;
assign W_R_STAGE_LUT[559] = 16'd168;
assign W_I_STAGE_LUT[559] = -16'd194;
assign W_R_STAGE_LUT[560] = 16'd167;
assign W_I_STAGE_LUT[560] = -16'd194;
assign W_R_STAGE_LUT[561] = 16'd167;
assign W_I_STAGE_LUT[561] = -16'd194;
assign W_R_STAGE_LUT[562] = 16'd167;
assign W_I_STAGE_LUT[562] = -16'd194;
assign W_R_STAGE_LUT[563] = 16'd166;
assign W_I_STAGE_LUT[563] = -16'd195;
assign W_R_STAGE_LUT[564] = 16'd166;
assign W_I_STAGE_LUT[564] = -16'd195;
assign W_R_STAGE_LUT[565] = 16'd166;
assign W_I_STAGE_LUT[565] = -16'd195;
assign W_R_STAGE_LUT[566] = 16'd165;
assign W_I_STAGE_LUT[566] = -16'd195;
assign W_R_STAGE_LUT[567] = 16'd165;
assign W_I_STAGE_LUT[567] = -16'd196;
assign W_R_STAGE_LUT[568] = 16'd165;
assign W_I_STAGE_LUT[568] = -16'd196;
assign W_R_STAGE_LUT[569] = 16'd165;
assign W_I_STAGE_LUT[569] = -16'd196;
assign W_R_STAGE_LUT[570] = 16'd164;
assign W_I_STAGE_LUT[570] = -16'd196;
assign W_R_STAGE_LUT[571] = 16'd164;
assign W_I_STAGE_LUT[571] = -16'd197;
assign W_R_STAGE_LUT[572] = 16'd164;
assign W_I_STAGE_LUT[572] = -16'd197;
assign W_R_STAGE_LUT[573] = 16'd163;
assign W_I_STAGE_LUT[573] = -16'd197;
assign W_R_STAGE_LUT[574] = 16'd163;
assign W_I_STAGE_LUT[574] = -16'd197;
assign W_R_STAGE_LUT[575] = 16'd163;
assign W_I_STAGE_LUT[575] = -16'd198;
assign W_R_STAGE_LUT[576] = 16'd162;
assign W_I_STAGE_LUT[576] = -16'd198;
assign W_R_STAGE_LUT[577] = 16'd162;
assign W_I_STAGE_LUT[577] = -16'd198;
assign W_R_STAGE_LUT[578] = 16'd162;
assign W_I_STAGE_LUT[578] = -16'd198;
assign W_R_STAGE_LUT[579] = 16'd161;
assign W_I_STAGE_LUT[579] = -16'd199;
assign W_R_STAGE_LUT[580] = 16'd161;
assign W_I_STAGE_LUT[580] = -16'd199;
assign W_R_STAGE_LUT[581] = 16'd161;
assign W_I_STAGE_LUT[581] = -16'd199;
assign W_R_STAGE_LUT[582] = 16'd161;
assign W_I_STAGE_LUT[582] = -16'd199;
assign W_R_STAGE_LUT[583] = 16'd160;
assign W_I_STAGE_LUT[583] = -16'd200;
assign W_R_STAGE_LUT[584] = 16'd160;
assign W_I_STAGE_LUT[584] = -16'd200;
assign W_R_STAGE_LUT[585] = 16'd160;
assign W_I_STAGE_LUT[585] = -16'd200;
assign W_R_STAGE_LUT[586] = 16'd159;
assign W_I_STAGE_LUT[586] = -16'd200;
assign W_R_STAGE_LUT[587] = 16'd159;
assign W_I_STAGE_LUT[587] = -16'd201;
assign W_R_STAGE_LUT[588] = 16'd159;
assign W_I_STAGE_LUT[588] = -16'd201;
assign W_R_STAGE_LUT[589] = 16'd158;
assign W_I_STAGE_LUT[589] = -16'd201;
assign W_R_STAGE_LUT[590] = 16'd158;
assign W_I_STAGE_LUT[590] = -16'd201;
assign W_R_STAGE_LUT[591] = 16'd158;
assign W_I_STAGE_LUT[591] = -16'd202;
assign W_R_STAGE_LUT[592] = 16'd157;
assign W_I_STAGE_LUT[592] = -16'd202;
assign W_R_STAGE_LUT[593] = 16'd157;
assign W_I_STAGE_LUT[593] = -16'd202;
assign W_R_STAGE_LUT[594] = 16'd157;
assign W_I_STAGE_LUT[594] = -16'd202;
assign W_R_STAGE_LUT[595] = 16'd157;
assign W_I_STAGE_LUT[595] = -16'd203;
assign W_R_STAGE_LUT[596] = 16'd156;
assign W_I_STAGE_LUT[596] = -16'd203;
assign W_R_STAGE_LUT[597] = 16'd156;
assign W_I_STAGE_LUT[597] = -16'd203;
assign W_R_STAGE_LUT[598] = 16'd156;
assign W_I_STAGE_LUT[598] = -16'd203;
assign W_R_STAGE_LUT[599] = 16'd155;
assign W_I_STAGE_LUT[599] = -16'd203;
assign W_R_STAGE_LUT[600] = 16'd155;
assign W_I_STAGE_LUT[600] = -16'd204;
assign W_R_STAGE_LUT[601] = 16'd155;
assign W_I_STAGE_LUT[601] = -16'd204;
assign W_R_STAGE_LUT[602] = 16'd154;
assign W_I_STAGE_LUT[602] = -16'd204;
assign W_R_STAGE_LUT[603] = 16'd154;
assign W_I_STAGE_LUT[603] = -16'd204;
assign W_R_STAGE_LUT[604] = 16'd154;
assign W_I_STAGE_LUT[604] = -16'd205;
assign W_R_STAGE_LUT[605] = 16'd153;
assign W_I_STAGE_LUT[605] = -16'd205;
assign W_R_STAGE_LUT[606] = 16'd153;
assign W_I_STAGE_LUT[606] = -16'd205;
assign W_R_STAGE_LUT[607] = 16'd153;
assign W_I_STAGE_LUT[607] = -16'd205;
assign W_R_STAGE_LUT[608] = 16'd152;
assign W_I_STAGE_LUT[608] = -16'd206;
assign W_R_STAGE_LUT[609] = 16'd152;
assign W_I_STAGE_LUT[609] = -16'd206;
assign W_R_STAGE_LUT[610] = 16'd152;
assign W_I_STAGE_LUT[610] = -16'd206;
assign W_R_STAGE_LUT[611] = 16'd152;
assign W_I_STAGE_LUT[611] = -16'd206;
assign W_R_STAGE_LUT[612] = 16'd151;
assign W_I_STAGE_LUT[612] = -16'd207;
assign W_R_STAGE_LUT[613] = 16'd151;
assign W_I_STAGE_LUT[613] = -16'd207;
assign W_R_STAGE_LUT[614] = 16'd151;
assign W_I_STAGE_LUT[614] = -16'd207;
assign W_R_STAGE_LUT[615] = 16'd150;
assign W_I_STAGE_LUT[615] = -16'd207;
assign W_R_STAGE_LUT[616] = 16'd150;
assign W_I_STAGE_LUT[616] = -16'd207;
assign W_R_STAGE_LUT[617] = 16'd150;
assign W_I_STAGE_LUT[617] = -16'd208;
assign W_R_STAGE_LUT[618] = 16'd149;
assign W_I_STAGE_LUT[618] = -16'd208;
assign W_R_STAGE_LUT[619] = 16'd149;
assign W_I_STAGE_LUT[619] = -16'd208;
assign W_R_STAGE_LUT[620] = 16'd149;
assign W_I_STAGE_LUT[620] = -16'd208;
assign W_R_STAGE_LUT[621] = 16'd148;
assign W_I_STAGE_LUT[621] = -16'd209;
assign W_R_STAGE_LUT[622] = 16'd148;
assign W_I_STAGE_LUT[622] = -16'd209;
assign W_R_STAGE_LUT[623] = 16'd148;
assign W_I_STAGE_LUT[623] = -16'd209;
assign W_R_STAGE_LUT[624] = 16'd147;
assign W_I_STAGE_LUT[624] = -16'd209;
assign W_R_STAGE_LUT[625] = 16'd147;
assign W_I_STAGE_LUT[625] = -16'd210;
assign W_R_STAGE_LUT[626] = 16'd147;
assign W_I_STAGE_LUT[626] = -16'd210;
assign W_R_STAGE_LUT[627] = 16'd146;
assign W_I_STAGE_LUT[627] = -16'd210;
assign W_R_STAGE_LUT[628] = 16'd146;
assign W_I_STAGE_LUT[628] = -16'd210;
assign W_R_STAGE_LUT[629] = 16'd146;
assign W_I_STAGE_LUT[629] = -16'd210;
assign W_R_STAGE_LUT[630] = 16'd145;
assign W_I_STAGE_LUT[630] = -16'd211;
assign W_R_STAGE_LUT[631] = 16'd145;
assign W_I_STAGE_LUT[631] = -16'd211;
assign W_R_STAGE_LUT[632] = 16'd145;
assign W_I_STAGE_LUT[632] = -16'd211;
assign W_R_STAGE_LUT[633] = 16'd145;
assign W_I_STAGE_LUT[633] = -16'd211;
assign W_R_STAGE_LUT[634] = 16'd144;
assign W_I_STAGE_LUT[634] = -16'd212;
assign W_R_STAGE_LUT[635] = 16'd144;
assign W_I_STAGE_LUT[635] = -16'd212;
assign W_R_STAGE_LUT[636] = 16'd144;
assign W_I_STAGE_LUT[636] = -16'd212;
assign W_R_STAGE_LUT[637] = 16'd143;
assign W_I_STAGE_LUT[637] = -16'd212;
assign W_R_STAGE_LUT[638] = 16'd143;
assign W_I_STAGE_LUT[638] = -16'd212;
assign W_R_STAGE_LUT[639] = 16'd143;
assign W_I_STAGE_LUT[639] = -16'd213;
assign W_R_STAGE_LUT[640] = 16'd142;
assign W_I_STAGE_LUT[640] = -16'd213;
assign W_R_STAGE_LUT[641] = 16'd142;
assign W_I_STAGE_LUT[641] = -16'd213;
assign W_R_STAGE_LUT[642] = 16'd142;
assign W_I_STAGE_LUT[642] = -16'd213;
assign W_R_STAGE_LUT[643] = 16'd141;
assign W_I_STAGE_LUT[643] = -16'd214;
assign W_R_STAGE_LUT[644] = 16'd141;
assign W_I_STAGE_LUT[644] = -16'd214;
assign W_R_STAGE_LUT[645] = 16'd141;
assign W_I_STAGE_LUT[645] = -16'd214;
assign W_R_STAGE_LUT[646] = 16'd140;
assign W_I_STAGE_LUT[646] = -16'd214;
assign W_R_STAGE_LUT[647] = 16'd140;
assign W_I_STAGE_LUT[647] = -16'd214;
assign W_R_STAGE_LUT[648] = 16'd140;
assign W_I_STAGE_LUT[648] = -16'd215;
assign W_R_STAGE_LUT[649] = 16'd139;
assign W_I_STAGE_LUT[649] = -16'd215;
assign W_R_STAGE_LUT[650] = 16'd139;
assign W_I_STAGE_LUT[650] = -16'd215;
assign W_R_STAGE_LUT[651] = 16'd139;
assign W_I_STAGE_LUT[651] = -16'd215;
assign W_R_STAGE_LUT[652] = 16'd138;
assign W_I_STAGE_LUT[652] = -16'd215;
assign W_R_STAGE_LUT[653] = 16'd138;
assign W_I_STAGE_LUT[653] = -16'd216;
assign W_R_STAGE_LUT[654] = 16'd138;
assign W_I_STAGE_LUT[654] = -16'd216;
assign W_R_STAGE_LUT[655] = 16'd137;
assign W_I_STAGE_LUT[655] = -16'd216;
assign W_R_STAGE_LUT[656] = 16'd137;
assign W_I_STAGE_LUT[656] = -16'd216;
assign W_R_STAGE_LUT[657] = 16'd137;
assign W_I_STAGE_LUT[657] = -16'd216;
assign W_R_STAGE_LUT[658] = 16'd136;
assign W_I_STAGE_LUT[658] = -16'd217;
assign W_R_STAGE_LUT[659] = 16'd136;
assign W_I_STAGE_LUT[659] = -16'd217;
assign W_R_STAGE_LUT[660] = 16'd136;
assign W_I_STAGE_LUT[660] = -16'd217;
assign W_R_STAGE_LUT[661] = 16'd135;
assign W_I_STAGE_LUT[661] = -16'd217;
assign W_R_STAGE_LUT[662] = 16'd135;
assign W_I_STAGE_LUT[662] = -16'd218;
assign W_R_STAGE_LUT[663] = 16'd135;
assign W_I_STAGE_LUT[663] = -16'd218;
assign W_R_STAGE_LUT[664] = 16'd134;
assign W_I_STAGE_LUT[664] = -16'd218;
assign W_R_STAGE_LUT[665] = 16'd134;
assign W_I_STAGE_LUT[665] = -16'd218;
assign W_R_STAGE_LUT[666] = 16'd134;
assign W_I_STAGE_LUT[666] = -16'd218;
assign W_R_STAGE_LUT[667] = 16'd133;
assign W_I_STAGE_LUT[667] = -16'd219;
assign W_R_STAGE_LUT[668] = 16'd133;
assign W_I_STAGE_LUT[668] = -16'd219;
assign W_R_STAGE_LUT[669] = 16'd133;
assign W_I_STAGE_LUT[669] = -16'd219;
assign W_R_STAGE_LUT[670] = 16'd132;
assign W_I_STAGE_LUT[670] = -16'd219;
assign W_R_STAGE_LUT[671] = 16'd132;
assign W_I_STAGE_LUT[671] = -16'd219;
assign W_R_STAGE_LUT[672] = 16'd132;
assign W_I_STAGE_LUT[672] = -16'd220;
assign W_R_STAGE_LUT[673] = 16'd131;
assign W_I_STAGE_LUT[673] = -16'd220;
assign W_R_STAGE_LUT[674] = 16'd131;
assign W_I_STAGE_LUT[674] = -16'd220;
assign W_R_STAGE_LUT[675] = 16'd131;
assign W_I_STAGE_LUT[675] = -16'd220;
assign W_R_STAGE_LUT[676] = 16'd130;
assign W_I_STAGE_LUT[676] = -16'd220;
assign W_R_STAGE_LUT[677] = 16'd130;
assign W_I_STAGE_LUT[677] = -16'd221;
assign W_R_STAGE_LUT[678] = 16'd130;
assign W_I_STAGE_LUT[678] = -16'd221;
assign W_R_STAGE_LUT[679] = 16'd129;
assign W_I_STAGE_LUT[679] = -16'd221;
assign W_R_STAGE_LUT[680] = 16'd129;
assign W_I_STAGE_LUT[680] = -16'd221;
assign W_R_STAGE_LUT[681] = 16'd129;
assign W_I_STAGE_LUT[681] = -16'd221;
assign W_R_STAGE_LUT[682] = 16'd128;
assign W_I_STAGE_LUT[682] = -16'd222;
assign W_R_STAGE_LUT[683] = 16'd128;
assign W_I_STAGE_LUT[683] = -16'd222;
assign W_R_STAGE_LUT[684] = 16'd128;
assign W_I_STAGE_LUT[684] = -16'd222;
assign W_R_STAGE_LUT[685] = 16'd127;
assign W_I_STAGE_LUT[685] = -16'd222;
assign W_R_STAGE_LUT[686] = 16'd127;
assign W_I_STAGE_LUT[686] = -16'd222;
assign W_R_STAGE_LUT[687] = 16'd127;
assign W_I_STAGE_LUT[687] = -16'd223;
assign W_R_STAGE_LUT[688] = 16'd126;
assign W_I_STAGE_LUT[688] = -16'd223;
assign W_R_STAGE_LUT[689] = 16'd126;
assign W_I_STAGE_LUT[689] = -16'd223;
assign W_R_STAGE_LUT[690] = 16'd125;
assign W_I_STAGE_LUT[690] = -16'd223;
assign W_R_STAGE_LUT[691] = 16'd125;
assign W_I_STAGE_LUT[691] = -16'd223;
assign W_R_STAGE_LUT[692] = 16'd125;
assign W_I_STAGE_LUT[692] = -16'd224;
assign W_R_STAGE_LUT[693] = 16'd124;
assign W_I_STAGE_LUT[693] = -16'd224;
assign W_R_STAGE_LUT[694] = 16'd124;
assign W_I_STAGE_LUT[694] = -16'd224;
assign W_R_STAGE_LUT[695] = 16'd124;
assign W_I_STAGE_LUT[695] = -16'd224;
assign W_R_STAGE_LUT[696] = 16'd123;
assign W_I_STAGE_LUT[696] = -16'd224;
assign W_R_STAGE_LUT[697] = 16'd123;
assign W_I_STAGE_LUT[697] = -16'd224;
assign W_R_STAGE_LUT[698] = 16'd123;
assign W_I_STAGE_LUT[698] = -16'd225;
assign W_R_STAGE_LUT[699] = 16'd122;
assign W_I_STAGE_LUT[699] = -16'd225;
assign W_R_STAGE_LUT[700] = 16'd122;
assign W_I_STAGE_LUT[700] = -16'd225;
assign W_R_STAGE_LUT[701] = 16'd122;
assign W_I_STAGE_LUT[701] = -16'd225;
assign W_R_STAGE_LUT[702] = 16'd121;
assign W_I_STAGE_LUT[702] = -16'd225;
assign W_R_STAGE_LUT[703] = 16'd121;
assign W_I_STAGE_LUT[703] = -16'd226;
assign W_R_STAGE_LUT[704] = 16'd121;
assign W_I_STAGE_LUT[704] = -16'd226;
assign W_R_STAGE_LUT[705] = 16'd120;
assign W_I_STAGE_LUT[705] = -16'd226;
assign W_R_STAGE_LUT[706] = 16'd120;
assign W_I_STAGE_LUT[706] = -16'd226;
assign W_R_STAGE_LUT[707] = 16'd120;
assign W_I_STAGE_LUT[707] = -16'd226;
assign W_R_STAGE_LUT[708] = 16'd119;
assign W_I_STAGE_LUT[708] = -16'd227;
assign W_R_STAGE_LUT[709] = 16'd119;
assign W_I_STAGE_LUT[709] = -16'd227;
assign W_R_STAGE_LUT[710] = 16'd119;
assign W_I_STAGE_LUT[710] = -16'd227;
assign W_R_STAGE_LUT[711] = 16'd118;
assign W_I_STAGE_LUT[711] = -16'd227;
assign W_R_STAGE_LUT[712] = 16'd118;
assign W_I_STAGE_LUT[712] = -16'd227;
assign W_R_STAGE_LUT[713] = 16'd118;
assign W_I_STAGE_LUT[713] = -16'd227;
assign W_R_STAGE_LUT[714] = 16'd117;
assign W_I_STAGE_LUT[714] = -16'd228;
assign W_R_STAGE_LUT[715] = 16'd117;
assign W_I_STAGE_LUT[715] = -16'd228;
assign W_R_STAGE_LUT[716] = 16'd117;
assign W_I_STAGE_LUT[716] = -16'd228;
assign W_R_STAGE_LUT[717] = 16'd116;
assign W_I_STAGE_LUT[717] = -16'd228;
assign W_R_STAGE_LUT[718] = 16'd116;
assign W_I_STAGE_LUT[718] = -16'd228;
assign W_R_STAGE_LUT[719] = 16'd115;
assign W_I_STAGE_LUT[719] = -16'd228;
assign W_R_STAGE_LUT[720] = 16'd115;
assign W_I_STAGE_LUT[720] = -16'd229;
assign W_R_STAGE_LUT[721] = 16'd115;
assign W_I_STAGE_LUT[721] = -16'd229;
assign W_R_STAGE_LUT[722] = 16'd114;
assign W_I_STAGE_LUT[722] = -16'd229;
assign W_R_STAGE_LUT[723] = 16'd114;
assign W_I_STAGE_LUT[723] = -16'd229;
assign W_R_STAGE_LUT[724] = 16'd114;
assign W_I_STAGE_LUT[724] = -16'd229;
assign W_R_STAGE_LUT[725] = 16'd113;
assign W_I_STAGE_LUT[725] = -16'd230;
assign W_R_STAGE_LUT[726] = 16'd113;
assign W_I_STAGE_LUT[726] = -16'd230;
assign W_R_STAGE_LUT[727] = 16'd113;
assign W_I_STAGE_LUT[727] = -16'd230;
assign W_R_STAGE_LUT[728] = 16'd112;
assign W_I_STAGE_LUT[728] = -16'd230;
assign W_R_STAGE_LUT[729] = 16'd112;
assign W_I_STAGE_LUT[729] = -16'd230;
assign W_R_STAGE_LUT[730] = 16'd112;
assign W_I_STAGE_LUT[730] = -16'd230;
assign W_R_STAGE_LUT[731] = 16'd111;
assign W_I_STAGE_LUT[731] = -16'd231;
assign W_R_STAGE_LUT[732] = 16'd111;
assign W_I_STAGE_LUT[732] = -16'd231;
assign W_R_STAGE_LUT[733] = 16'd111;
assign W_I_STAGE_LUT[733] = -16'd231;
assign W_R_STAGE_LUT[734] = 16'd110;
assign W_I_STAGE_LUT[734] = -16'd231;
assign W_R_STAGE_LUT[735] = 16'd110;
assign W_I_STAGE_LUT[735] = -16'd231;
assign W_R_STAGE_LUT[736] = 16'd109;
assign W_I_STAGE_LUT[736] = -16'd231;
assign W_R_STAGE_LUT[737] = 16'd109;
assign W_I_STAGE_LUT[737] = -16'd232;
assign W_R_STAGE_LUT[738] = 16'd109;
assign W_I_STAGE_LUT[738] = -16'd232;
assign W_R_STAGE_LUT[739] = 16'd108;
assign W_I_STAGE_LUT[739] = -16'd232;
assign W_R_STAGE_LUT[740] = 16'd108;
assign W_I_STAGE_LUT[740] = -16'd232;
assign W_R_STAGE_LUT[741] = 16'd108;
assign W_I_STAGE_LUT[741] = -16'd232;
assign W_R_STAGE_LUT[742] = 16'd107;
assign W_I_STAGE_LUT[742] = -16'd232;
assign W_R_STAGE_LUT[743] = 16'd107;
assign W_I_STAGE_LUT[743] = -16'd233;
assign W_R_STAGE_LUT[744] = 16'd107;
assign W_I_STAGE_LUT[744] = -16'd233;
assign W_R_STAGE_LUT[745] = 16'd106;
assign W_I_STAGE_LUT[745] = -16'd233;
assign W_R_STAGE_LUT[746] = 16'd106;
assign W_I_STAGE_LUT[746] = -16'd233;
assign W_R_STAGE_LUT[747] = 16'd106;
assign W_I_STAGE_LUT[747] = -16'd233;
assign W_R_STAGE_LUT[748] = 16'd105;
assign W_I_STAGE_LUT[748] = -16'd233;
assign W_R_STAGE_LUT[749] = 16'd105;
assign W_I_STAGE_LUT[749] = -16'd234;
assign W_R_STAGE_LUT[750] = 16'd104;
assign W_I_STAGE_LUT[750] = -16'd234;
assign W_R_STAGE_LUT[751] = 16'd104;
assign W_I_STAGE_LUT[751] = -16'd234;
assign W_R_STAGE_LUT[752] = 16'd104;
assign W_I_STAGE_LUT[752] = -16'd234;
assign W_R_STAGE_LUT[753] = 16'd103;
assign W_I_STAGE_LUT[753] = -16'd234;
assign W_R_STAGE_LUT[754] = 16'd103;
assign W_I_STAGE_LUT[754] = -16'd234;
assign W_R_STAGE_LUT[755] = 16'd103;
assign W_I_STAGE_LUT[755] = -16'd235;
assign W_R_STAGE_LUT[756] = 16'd102;
assign W_I_STAGE_LUT[756] = -16'd235;
assign W_R_STAGE_LUT[757] = 16'd102;
assign W_I_STAGE_LUT[757] = -16'd235;
assign W_R_STAGE_LUT[758] = 16'd102;
assign W_I_STAGE_LUT[758] = -16'd235;
assign W_R_STAGE_LUT[759] = 16'd101;
assign W_I_STAGE_LUT[759] = -16'd235;
assign W_R_STAGE_LUT[760] = 16'd101;
assign W_I_STAGE_LUT[760] = -16'd235;
assign W_R_STAGE_LUT[761] = 16'd101;
assign W_I_STAGE_LUT[761] = -16'd235;
assign W_R_STAGE_LUT[762] = 16'd100;
assign W_I_STAGE_LUT[762] = -16'd236;
assign W_R_STAGE_LUT[763] = 16'd100;
assign W_I_STAGE_LUT[763] = -16'd236;
assign W_R_STAGE_LUT[764] = 16'd99;
assign W_I_STAGE_LUT[764] = -16'd236;
assign W_R_STAGE_LUT[765] = 16'd99;
assign W_I_STAGE_LUT[765] = -16'd236;
assign W_R_STAGE_LUT[766] = 16'd99;
assign W_I_STAGE_LUT[766] = -16'd236;
assign W_R_STAGE_LUT[767] = 16'd98;
assign W_I_STAGE_LUT[767] = -16'd236;
assign W_R_STAGE_LUT[768] = 16'd98;
assign W_I_STAGE_LUT[768] = -16'd237;
assign W_R_STAGE_LUT[769] = 16'd98;
assign W_I_STAGE_LUT[769] = -16'd237;
assign W_R_STAGE_LUT[770] = 16'd97;
assign W_I_STAGE_LUT[770] = -16'd237;
assign W_R_STAGE_LUT[771] = 16'd97;
assign W_I_STAGE_LUT[771] = -16'd237;
assign W_R_STAGE_LUT[772] = 16'd97;
assign W_I_STAGE_LUT[772] = -16'd237;
assign W_R_STAGE_LUT[773] = 16'd96;
assign W_I_STAGE_LUT[773] = -16'd237;
assign W_R_STAGE_LUT[774] = 16'd96;
assign W_I_STAGE_LUT[774] = -16'd237;
assign W_R_STAGE_LUT[775] = 16'd95;
assign W_I_STAGE_LUT[775] = -16'd238;
assign W_R_STAGE_LUT[776] = 16'd95;
assign W_I_STAGE_LUT[776] = -16'd238;
assign W_R_STAGE_LUT[777] = 16'd95;
assign W_I_STAGE_LUT[777] = -16'd238;
assign W_R_STAGE_LUT[778] = 16'd94;
assign W_I_STAGE_LUT[778] = -16'd238;
assign W_R_STAGE_LUT[779] = 16'd94;
assign W_I_STAGE_LUT[779] = -16'd238;
assign W_R_STAGE_LUT[780] = 16'd94;
assign W_I_STAGE_LUT[780] = -16'd238;
assign W_R_STAGE_LUT[781] = 16'd93;
assign W_I_STAGE_LUT[781] = -16'd238;
assign W_R_STAGE_LUT[782] = 16'd93;
assign W_I_STAGE_LUT[782] = -16'd239;
assign W_R_STAGE_LUT[783] = 16'd92;
assign W_I_STAGE_LUT[783] = -16'd239;
assign W_R_STAGE_LUT[784] = 16'd92;
assign W_I_STAGE_LUT[784] = -16'd239;
assign W_R_STAGE_LUT[785] = 16'd92;
assign W_I_STAGE_LUT[785] = -16'd239;
assign W_R_STAGE_LUT[786] = 16'd91;
assign W_I_STAGE_LUT[786] = -16'd239;
assign W_R_STAGE_LUT[787] = 16'd91;
assign W_I_STAGE_LUT[787] = -16'd239;
assign W_R_STAGE_LUT[788] = 16'd91;
assign W_I_STAGE_LUT[788] = -16'd239;
assign W_R_STAGE_LUT[789] = 16'd90;
assign W_I_STAGE_LUT[789] = -16'd240;
assign W_R_STAGE_LUT[790] = 16'd90;
assign W_I_STAGE_LUT[790] = -16'd240;
assign W_R_STAGE_LUT[791] = 16'd90;
assign W_I_STAGE_LUT[791] = -16'd240;
assign W_R_STAGE_LUT[792] = 16'd89;
assign W_I_STAGE_LUT[792] = -16'd240;
assign W_R_STAGE_LUT[793] = 16'd89;
assign W_I_STAGE_LUT[793] = -16'd240;
assign W_R_STAGE_LUT[794] = 16'd88;
assign W_I_STAGE_LUT[794] = -16'd240;
assign W_R_STAGE_LUT[795] = 16'd88;
assign W_I_STAGE_LUT[795] = -16'd240;
assign W_R_STAGE_LUT[796] = 16'd88;
assign W_I_STAGE_LUT[796] = -16'd241;
assign W_R_STAGE_LUT[797] = 16'd87;
assign W_I_STAGE_LUT[797] = -16'd241;
assign W_R_STAGE_LUT[798] = 16'd87;
assign W_I_STAGE_LUT[798] = -16'd241;
assign W_R_STAGE_LUT[799] = 16'd87;
assign W_I_STAGE_LUT[799] = -16'd241;
assign W_R_STAGE_LUT[800] = 16'd86;
assign W_I_STAGE_LUT[800] = -16'd241;
assign W_R_STAGE_LUT[801] = 16'd86;
assign W_I_STAGE_LUT[801] = -16'd241;
assign W_R_STAGE_LUT[802] = 16'd86;
assign W_I_STAGE_LUT[802] = -16'd241;
assign W_R_STAGE_LUT[803] = 16'd85;
assign W_I_STAGE_LUT[803] = -16'd241;
assign W_R_STAGE_LUT[804] = 16'd85;
assign W_I_STAGE_LUT[804] = -16'd242;
assign W_R_STAGE_LUT[805] = 16'd84;
assign W_I_STAGE_LUT[805] = -16'd242;
assign W_R_STAGE_LUT[806] = 16'd84;
assign W_I_STAGE_LUT[806] = -16'd242;
assign W_R_STAGE_LUT[807] = 16'd84;
assign W_I_STAGE_LUT[807] = -16'd242;
assign W_R_STAGE_LUT[808] = 16'd83;
assign W_I_STAGE_LUT[808] = -16'd242;
assign W_R_STAGE_LUT[809] = 16'd83;
assign W_I_STAGE_LUT[809] = -16'd242;
assign W_R_STAGE_LUT[810] = 16'd83;
assign W_I_STAGE_LUT[810] = -16'd242;
assign W_R_STAGE_LUT[811] = 16'd82;
assign W_I_STAGE_LUT[811] = -16'd242;
assign W_R_STAGE_LUT[812] = 16'd82;
assign W_I_STAGE_LUT[812] = -16'd243;
assign W_R_STAGE_LUT[813] = 16'd81;
assign W_I_STAGE_LUT[813] = -16'd243;
assign W_R_STAGE_LUT[814] = 16'd81;
assign W_I_STAGE_LUT[814] = -16'd243;
assign W_R_STAGE_LUT[815] = 16'd81;
assign W_I_STAGE_LUT[815] = -16'd243;
assign W_R_STAGE_LUT[816] = 16'd80;
assign W_I_STAGE_LUT[816] = -16'd243;
assign W_R_STAGE_LUT[817] = 16'd80;
assign W_I_STAGE_LUT[817] = -16'd243;
assign W_R_STAGE_LUT[818] = 16'd80;
assign W_I_STAGE_LUT[818] = -16'd243;
assign W_R_STAGE_LUT[819] = 16'd79;
assign W_I_STAGE_LUT[819] = -16'd243;
assign W_R_STAGE_LUT[820] = 16'd79;
assign W_I_STAGE_LUT[820] = -16'd244;
assign W_R_STAGE_LUT[821] = 16'd78;
assign W_I_STAGE_LUT[821] = -16'd244;
assign W_R_STAGE_LUT[822] = 16'd78;
assign W_I_STAGE_LUT[822] = -16'd244;
assign W_R_STAGE_LUT[823] = 16'd78;
assign W_I_STAGE_LUT[823] = -16'd244;
assign W_R_STAGE_LUT[824] = 16'd77;
assign W_I_STAGE_LUT[824] = -16'd244;
assign W_R_STAGE_LUT[825] = 16'd77;
assign W_I_STAGE_LUT[825] = -16'd244;
assign W_R_STAGE_LUT[826] = 16'd77;
assign W_I_STAGE_LUT[826] = -16'd244;
assign W_R_STAGE_LUT[827] = 16'd76;
assign W_I_STAGE_LUT[827] = -16'd244;
assign W_R_STAGE_LUT[828] = 16'd76;
assign W_I_STAGE_LUT[828] = -16'd245;
assign W_R_STAGE_LUT[829] = 16'd75;
assign W_I_STAGE_LUT[829] = -16'd245;
assign W_R_STAGE_LUT[830] = 16'd75;
assign W_I_STAGE_LUT[830] = -16'd245;
assign W_R_STAGE_LUT[831] = 16'd75;
assign W_I_STAGE_LUT[831] = -16'd245;
assign W_R_STAGE_LUT[832] = 16'd74;
assign W_I_STAGE_LUT[832] = -16'd245;
assign W_R_STAGE_LUT[833] = 16'd74;
assign W_I_STAGE_LUT[833] = -16'd245;
assign W_R_STAGE_LUT[834] = 16'd74;
assign W_I_STAGE_LUT[834] = -16'd245;
assign W_R_STAGE_LUT[835] = 16'd73;
assign W_I_STAGE_LUT[835] = -16'd245;
assign W_R_STAGE_LUT[836] = 16'd73;
assign W_I_STAGE_LUT[836] = -16'd245;
assign W_R_STAGE_LUT[837] = 16'd72;
assign W_I_STAGE_LUT[837] = -16'd246;
assign W_R_STAGE_LUT[838] = 16'd72;
assign W_I_STAGE_LUT[838] = -16'd246;
assign W_R_STAGE_LUT[839] = 16'd72;
assign W_I_STAGE_LUT[839] = -16'd246;
assign W_R_STAGE_LUT[840] = 16'd71;
assign W_I_STAGE_LUT[840] = -16'd246;
assign W_R_STAGE_LUT[841] = 16'd71;
assign W_I_STAGE_LUT[841] = -16'd246;
assign W_R_STAGE_LUT[842] = 16'd71;
assign W_I_STAGE_LUT[842] = -16'd246;
assign W_R_STAGE_LUT[843] = 16'd70;
assign W_I_STAGE_LUT[843] = -16'd246;
assign W_R_STAGE_LUT[844] = 16'd70;
assign W_I_STAGE_LUT[844] = -16'd246;
assign W_R_STAGE_LUT[845] = 16'd69;
assign W_I_STAGE_LUT[845] = -16'd246;
assign W_R_STAGE_LUT[846] = 16'd69;
assign W_I_STAGE_LUT[846] = -16'd247;
assign W_R_STAGE_LUT[847] = 16'd69;
assign W_I_STAGE_LUT[847] = -16'd247;
assign W_R_STAGE_LUT[848] = 16'd68;
assign W_I_STAGE_LUT[848] = -16'd247;
assign W_R_STAGE_LUT[849] = 16'd68;
assign W_I_STAGE_LUT[849] = -16'd247;
assign W_R_STAGE_LUT[850] = 16'd68;
assign W_I_STAGE_LUT[850] = -16'd247;
assign W_R_STAGE_LUT[851] = 16'd67;
assign W_I_STAGE_LUT[851] = -16'd247;
assign W_R_STAGE_LUT[852] = 16'd67;
assign W_I_STAGE_LUT[852] = -16'd247;
assign W_R_STAGE_LUT[853] = 16'd66;
assign W_I_STAGE_LUT[853] = -16'd247;
assign W_R_STAGE_LUT[854] = 16'd66;
assign W_I_STAGE_LUT[854] = -16'd247;
assign W_R_STAGE_LUT[855] = 16'd66;
assign W_I_STAGE_LUT[855] = -16'd247;
assign W_R_STAGE_LUT[856] = 16'd65;
assign W_I_STAGE_LUT[856] = -16'd248;
assign W_R_STAGE_LUT[857] = 16'd65;
assign W_I_STAGE_LUT[857] = -16'd248;
assign W_R_STAGE_LUT[858] = 16'd64;
assign W_I_STAGE_LUT[858] = -16'd248;
assign W_R_STAGE_LUT[859] = 16'd64;
assign W_I_STAGE_LUT[859] = -16'd248;
assign W_R_STAGE_LUT[860] = 16'd64;
assign W_I_STAGE_LUT[860] = -16'd248;
assign W_R_STAGE_LUT[861] = 16'd63;
assign W_I_STAGE_LUT[861] = -16'd248;
assign W_R_STAGE_LUT[862] = 16'd63;
assign W_I_STAGE_LUT[862] = -16'd248;
assign W_R_STAGE_LUT[863] = 16'd63;
assign W_I_STAGE_LUT[863] = -16'd248;
assign W_R_STAGE_LUT[864] = 16'd62;
assign W_I_STAGE_LUT[864] = -16'd248;
assign W_R_STAGE_LUT[865] = 16'd62;
assign W_I_STAGE_LUT[865] = -16'd248;
assign W_R_STAGE_LUT[866] = 16'd61;
assign W_I_STAGE_LUT[866] = -16'd249;
assign W_R_STAGE_LUT[867] = 16'd61;
assign W_I_STAGE_LUT[867] = -16'd249;
assign W_R_STAGE_LUT[868] = 16'd61;
assign W_I_STAGE_LUT[868] = -16'd249;
assign W_R_STAGE_LUT[869] = 16'd60;
assign W_I_STAGE_LUT[869] = -16'd249;
assign W_R_STAGE_LUT[870] = 16'd60;
assign W_I_STAGE_LUT[870] = -16'd249;
assign W_R_STAGE_LUT[871] = 16'd60;
assign W_I_STAGE_LUT[871] = -16'd249;
assign W_R_STAGE_LUT[872] = 16'd59;
assign W_I_STAGE_LUT[872] = -16'd249;
assign W_R_STAGE_LUT[873] = 16'd59;
assign W_I_STAGE_LUT[873] = -16'd249;
assign W_R_STAGE_LUT[874] = 16'd58;
assign W_I_STAGE_LUT[874] = -16'd249;
assign W_R_STAGE_LUT[875] = 16'd58;
assign W_I_STAGE_LUT[875] = -16'd249;
assign W_R_STAGE_LUT[876] = 16'd58;
assign W_I_STAGE_LUT[876] = -16'd249;
assign W_R_STAGE_LUT[877] = 16'd57;
assign W_I_STAGE_LUT[877] = -16'd250;
assign W_R_STAGE_LUT[878] = 16'd57;
assign W_I_STAGE_LUT[878] = -16'd250;
assign W_R_STAGE_LUT[879] = 16'd56;
assign W_I_STAGE_LUT[879] = -16'd250;
assign W_R_STAGE_LUT[880] = 16'd56;
assign W_I_STAGE_LUT[880] = -16'd250;
assign W_R_STAGE_LUT[881] = 16'd56;
assign W_I_STAGE_LUT[881] = -16'd250;
assign W_R_STAGE_LUT[882] = 16'd55;
assign W_I_STAGE_LUT[882] = -16'd250;
assign W_R_STAGE_LUT[883] = 16'd55;
assign W_I_STAGE_LUT[883] = -16'd250;
assign W_R_STAGE_LUT[884] = 16'd55;
assign W_I_STAGE_LUT[884] = -16'd250;
assign W_R_STAGE_LUT[885] = 16'd54;
assign W_I_STAGE_LUT[885] = -16'd250;
assign W_R_STAGE_LUT[886] = 16'd54;
assign W_I_STAGE_LUT[886] = -16'd250;
assign W_R_STAGE_LUT[887] = 16'd53;
assign W_I_STAGE_LUT[887] = -16'd250;
assign W_R_STAGE_LUT[888] = 16'd53;
assign W_I_STAGE_LUT[888] = -16'd250;
assign W_R_STAGE_LUT[889] = 16'd53;
assign W_I_STAGE_LUT[889] = -16'd251;
assign W_R_STAGE_LUT[890] = 16'd52;
assign W_I_STAGE_LUT[890] = -16'd251;
assign W_R_STAGE_LUT[891] = 16'd52;
assign W_I_STAGE_LUT[891] = -16'd251;
assign W_R_STAGE_LUT[892] = 16'd51;
assign W_I_STAGE_LUT[892] = -16'd251;
assign W_R_STAGE_LUT[893] = 16'd51;
assign W_I_STAGE_LUT[893] = -16'd251;
assign W_R_STAGE_LUT[894] = 16'd51;
assign W_I_STAGE_LUT[894] = -16'd251;
assign W_R_STAGE_LUT[895] = 16'd50;
assign W_I_STAGE_LUT[895] = -16'd251;
assign W_R_STAGE_LUT[896] = 16'd50;
assign W_I_STAGE_LUT[896] = -16'd251;
assign W_R_STAGE_LUT[897] = 16'd50;
assign W_I_STAGE_LUT[897] = -16'd251;
assign W_R_STAGE_LUT[898] = 16'd49;
assign W_I_STAGE_LUT[898] = -16'd251;
assign W_R_STAGE_LUT[899] = 16'd49;
assign W_I_STAGE_LUT[899] = -16'd251;
assign W_R_STAGE_LUT[900] = 16'd48;
assign W_I_STAGE_LUT[900] = -16'd251;
assign W_R_STAGE_LUT[901] = 16'd48;
assign W_I_STAGE_LUT[901] = -16'd251;
assign W_R_STAGE_LUT[902] = 16'd48;
assign W_I_STAGE_LUT[902] = -16'd252;
assign W_R_STAGE_LUT[903] = 16'd47;
assign W_I_STAGE_LUT[903] = -16'd252;
assign W_R_STAGE_LUT[904] = 16'd47;
assign W_I_STAGE_LUT[904] = -16'd252;
assign W_R_STAGE_LUT[905] = 16'd46;
assign W_I_STAGE_LUT[905] = -16'd252;
assign W_R_STAGE_LUT[906] = 16'd46;
assign W_I_STAGE_LUT[906] = -16'd252;
assign W_R_STAGE_LUT[907] = 16'd46;
assign W_I_STAGE_LUT[907] = -16'd252;
assign W_R_STAGE_LUT[908] = 16'd45;
assign W_I_STAGE_LUT[908] = -16'd252;
assign W_R_STAGE_LUT[909] = 16'd45;
assign W_I_STAGE_LUT[909] = -16'd252;
assign W_R_STAGE_LUT[910] = 16'd45;
assign W_I_STAGE_LUT[910] = -16'd252;
assign W_R_STAGE_LUT[911] = 16'd44;
assign W_I_STAGE_LUT[911] = -16'd252;
assign W_R_STAGE_LUT[912] = 16'd44;
assign W_I_STAGE_LUT[912] = -16'd252;
assign W_R_STAGE_LUT[913] = 16'd43;
assign W_I_STAGE_LUT[913] = -16'd252;
assign W_R_STAGE_LUT[914] = 16'd43;
assign W_I_STAGE_LUT[914] = -16'd252;
assign W_R_STAGE_LUT[915] = 16'd43;
assign W_I_STAGE_LUT[915] = -16'd252;
assign W_R_STAGE_LUT[916] = 16'd42;
assign W_I_STAGE_LUT[916] = -16'd252;
assign W_R_STAGE_LUT[917] = 16'd42;
assign W_I_STAGE_LUT[917] = -16'd253;
assign W_R_STAGE_LUT[918] = 16'd41;
assign W_I_STAGE_LUT[918] = -16'd253;
assign W_R_STAGE_LUT[919] = 16'd41;
assign W_I_STAGE_LUT[919] = -16'd253;
assign W_R_STAGE_LUT[920] = 16'd41;
assign W_I_STAGE_LUT[920] = -16'd253;
assign W_R_STAGE_LUT[921] = 16'd40;
assign W_I_STAGE_LUT[921] = -16'd253;
assign W_R_STAGE_LUT[922] = 16'd40;
assign W_I_STAGE_LUT[922] = -16'd253;
assign W_R_STAGE_LUT[923] = 16'd40;
assign W_I_STAGE_LUT[923] = -16'd253;
assign W_R_STAGE_LUT[924] = 16'd39;
assign W_I_STAGE_LUT[924] = -16'd253;
assign W_R_STAGE_LUT[925] = 16'd39;
assign W_I_STAGE_LUT[925] = -16'd253;
assign W_R_STAGE_LUT[926] = 16'd38;
assign W_I_STAGE_LUT[926] = -16'd253;
assign W_R_STAGE_LUT[927] = 16'd38;
assign W_I_STAGE_LUT[927] = -16'd253;
assign W_R_STAGE_LUT[928] = 16'd38;
assign W_I_STAGE_LUT[928] = -16'd253;
assign W_R_STAGE_LUT[929] = 16'd37;
assign W_I_STAGE_LUT[929] = -16'd253;
assign W_R_STAGE_LUT[930] = 16'd37;
assign W_I_STAGE_LUT[930] = -16'd253;
assign W_R_STAGE_LUT[931] = 16'd36;
assign W_I_STAGE_LUT[931] = -16'd253;
assign W_R_STAGE_LUT[932] = 16'd36;
assign W_I_STAGE_LUT[932] = -16'd253;
assign W_R_STAGE_LUT[933] = 16'd36;
assign W_I_STAGE_LUT[933] = -16'd254;
assign W_R_STAGE_LUT[934] = 16'd35;
assign W_I_STAGE_LUT[934] = -16'd254;
assign W_R_STAGE_LUT[935] = 16'd35;
assign W_I_STAGE_LUT[935] = -16'd254;
assign W_R_STAGE_LUT[936] = 16'd34;
assign W_I_STAGE_LUT[936] = -16'd254;
assign W_R_STAGE_LUT[937] = 16'd34;
assign W_I_STAGE_LUT[937] = -16'd254;
assign W_R_STAGE_LUT[938] = 16'd34;
assign W_I_STAGE_LUT[938] = -16'd254;
assign W_R_STAGE_LUT[939] = 16'd33;
assign W_I_STAGE_LUT[939] = -16'd254;
assign W_R_STAGE_LUT[940] = 16'd33;
assign W_I_STAGE_LUT[940] = -16'd254;
assign W_R_STAGE_LUT[941] = 16'd33;
assign W_I_STAGE_LUT[941] = -16'd254;
assign W_R_STAGE_LUT[942] = 16'd32;
assign W_I_STAGE_LUT[942] = -16'd254;
assign W_R_STAGE_LUT[943] = 16'd32;
assign W_I_STAGE_LUT[943] = -16'd254;
assign W_R_STAGE_LUT[944] = 16'd31;
assign W_I_STAGE_LUT[944] = -16'd254;
assign W_R_STAGE_LUT[945] = 16'd31;
assign W_I_STAGE_LUT[945] = -16'd254;
assign W_R_STAGE_LUT[946] = 16'd31;
assign W_I_STAGE_LUT[946] = -16'd254;
assign W_R_STAGE_LUT[947] = 16'd30;
assign W_I_STAGE_LUT[947] = -16'd254;
assign W_R_STAGE_LUT[948] = 16'd30;
assign W_I_STAGE_LUT[948] = -16'd254;
assign W_R_STAGE_LUT[949] = 16'd29;
assign W_I_STAGE_LUT[949] = -16'd254;
assign W_R_STAGE_LUT[950] = 16'd29;
assign W_I_STAGE_LUT[950] = -16'd254;
assign W_R_STAGE_LUT[951] = 16'd29;
assign W_I_STAGE_LUT[951] = -16'd254;
assign W_R_STAGE_LUT[952] = 16'd28;
assign W_I_STAGE_LUT[952] = -16'd254;
assign W_R_STAGE_LUT[953] = 16'd28;
assign W_I_STAGE_LUT[953] = -16'd254;
assign W_R_STAGE_LUT[954] = 16'd27;
assign W_I_STAGE_LUT[954] = -16'd255;
assign W_R_STAGE_LUT[955] = 16'd27;
assign W_I_STAGE_LUT[955] = -16'd255;
assign W_R_STAGE_LUT[956] = 16'd27;
assign W_I_STAGE_LUT[956] = -16'd255;
assign W_R_STAGE_LUT[957] = 16'd26;
assign W_I_STAGE_LUT[957] = -16'd255;
assign W_R_STAGE_LUT[958] = 16'd26;
assign W_I_STAGE_LUT[958] = -16'd255;
assign W_R_STAGE_LUT[959] = 16'd25;
assign W_I_STAGE_LUT[959] = -16'd255;
assign W_R_STAGE_LUT[960] = 16'd25;
assign W_I_STAGE_LUT[960] = -16'd255;
assign W_R_STAGE_LUT[961] = 16'd25;
assign W_I_STAGE_LUT[961] = -16'd255;
assign W_R_STAGE_LUT[962] = 16'd24;
assign W_I_STAGE_LUT[962] = -16'd255;
assign W_R_STAGE_LUT[963] = 16'd24;
assign W_I_STAGE_LUT[963] = -16'd255;
assign W_R_STAGE_LUT[964] = 16'd24;
assign W_I_STAGE_LUT[964] = -16'd255;
assign W_R_STAGE_LUT[965] = 16'd23;
assign W_I_STAGE_LUT[965] = -16'd255;
assign W_R_STAGE_LUT[966] = 16'd23;
assign W_I_STAGE_LUT[966] = -16'd255;
assign W_R_STAGE_LUT[967] = 16'd22;
assign W_I_STAGE_LUT[967] = -16'd255;
assign W_R_STAGE_LUT[968] = 16'd22;
assign W_I_STAGE_LUT[968] = -16'd255;
assign W_R_STAGE_LUT[969] = 16'd22;
assign W_I_STAGE_LUT[969] = -16'd255;
assign W_R_STAGE_LUT[970] = 16'd21;
assign W_I_STAGE_LUT[970] = -16'd255;
assign W_R_STAGE_LUT[971] = 16'd21;
assign W_I_STAGE_LUT[971] = -16'd255;
assign W_R_STAGE_LUT[972] = 16'd20;
assign W_I_STAGE_LUT[972] = -16'd255;
assign W_R_STAGE_LUT[973] = 16'd20;
assign W_I_STAGE_LUT[973] = -16'd255;
assign W_R_STAGE_LUT[974] = 16'd20;
assign W_I_STAGE_LUT[974] = -16'd255;
assign W_R_STAGE_LUT[975] = 16'd19;
assign W_I_STAGE_LUT[975] = -16'd255;
assign W_R_STAGE_LUT[976] = 16'd19;
assign W_I_STAGE_LUT[976] = -16'd255;
assign W_R_STAGE_LUT[977] = 16'd18;
assign W_I_STAGE_LUT[977] = -16'd255;
assign W_R_STAGE_LUT[978] = 16'd18;
assign W_I_STAGE_LUT[978] = -16'd255;
assign W_R_STAGE_LUT[979] = 16'd18;
assign W_I_STAGE_LUT[979] = -16'd255;
assign W_R_STAGE_LUT[980] = 16'd17;
assign W_I_STAGE_LUT[980] = -16'd255;
assign W_R_STAGE_LUT[981] = 16'd17;
assign W_I_STAGE_LUT[981] = -16'd255;
assign W_R_STAGE_LUT[982] = 16'd16;
assign W_I_STAGE_LUT[982] = -16'd255;
assign W_R_STAGE_LUT[983] = 16'd16;
assign W_I_STAGE_LUT[983] = -16'd255;
assign W_R_STAGE_LUT[984] = 16'd16;
assign W_I_STAGE_LUT[984] = -16'd256;
assign W_R_STAGE_LUT[985] = 16'd15;
assign W_I_STAGE_LUT[985] = -16'd256;
assign W_R_STAGE_LUT[986] = 16'd15;
assign W_I_STAGE_LUT[986] = -16'd256;
assign W_R_STAGE_LUT[987] = 16'd15;
assign W_I_STAGE_LUT[987] = -16'd256;
assign W_R_STAGE_LUT[988] = 16'd14;
assign W_I_STAGE_LUT[988] = -16'd256;
assign W_R_STAGE_LUT[989] = 16'd14;
assign W_I_STAGE_LUT[989] = -16'd256;
assign W_R_STAGE_LUT[990] = 16'd13;
assign W_I_STAGE_LUT[990] = -16'd256;
assign W_R_STAGE_LUT[991] = 16'd13;
assign W_I_STAGE_LUT[991] = -16'd256;
assign W_R_STAGE_LUT[992] = 16'd13;
assign W_I_STAGE_LUT[992] = -16'd256;
assign W_R_STAGE_LUT[993] = 16'd12;
assign W_I_STAGE_LUT[993] = -16'd256;
assign W_R_STAGE_LUT[994] = 16'd12;
assign W_I_STAGE_LUT[994] = -16'd256;
assign W_R_STAGE_LUT[995] = 16'd11;
assign W_I_STAGE_LUT[995] = -16'd256;
assign W_R_STAGE_LUT[996] = 16'd11;
assign W_I_STAGE_LUT[996] = -16'd256;
assign W_R_STAGE_LUT[997] = 16'd11;
assign W_I_STAGE_LUT[997] = -16'd256;
assign W_R_STAGE_LUT[998] = 16'd10;
assign W_I_STAGE_LUT[998] = -16'd256;
assign W_R_STAGE_LUT[999] = 16'd10;
assign W_I_STAGE_LUT[999] = -16'd256;
assign W_R_STAGE_LUT[1000] = 16'd9;
assign W_I_STAGE_LUT[1000] = -16'd256;
assign W_R_STAGE_LUT[1001] = 16'd9;
assign W_I_STAGE_LUT[1001] = -16'd256;
assign W_R_STAGE_LUT[1002] = 16'd9;
assign W_I_STAGE_LUT[1002] = -16'd256;
assign W_R_STAGE_LUT[1003] = 16'd8;
assign W_I_STAGE_LUT[1003] = -16'd256;
assign W_R_STAGE_LUT[1004] = 16'd8;
assign W_I_STAGE_LUT[1004] = -16'd256;
assign W_R_STAGE_LUT[1005] = 16'd7;
assign W_I_STAGE_LUT[1005] = -16'd256;
assign W_R_STAGE_LUT[1006] = 16'd7;
assign W_I_STAGE_LUT[1006] = -16'd256;
assign W_R_STAGE_LUT[1007] = 16'd7;
assign W_I_STAGE_LUT[1007] = -16'd256;
assign W_R_STAGE_LUT[1008] = 16'd6;
assign W_I_STAGE_LUT[1008] = -16'd256;
assign W_R_STAGE_LUT[1009] = 16'd6;
assign W_I_STAGE_LUT[1009] = -16'd256;
assign W_R_STAGE_LUT[1010] = 16'd5;
assign W_I_STAGE_LUT[1010] = -16'd256;
assign W_R_STAGE_LUT[1011] = 16'd5;
assign W_I_STAGE_LUT[1011] = -16'd256;
assign W_R_STAGE_LUT[1012] = 16'd5;
assign W_I_STAGE_LUT[1012] = -16'd256;
assign W_R_STAGE_LUT[1013] = 16'd4;
assign W_I_STAGE_LUT[1013] = -16'd256;
assign W_R_STAGE_LUT[1014] = 16'd4;
assign W_I_STAGE_LUT[1014] = -16'd256;
assign W_R_STAGE_LUT[1015] = 16'd4;
assign W_I_STAGE_LUT[1015] = -16'd256;
assign W_R_STAGE_LUT[1016] = 16'd3;
assign W_I_STAGE_LUT[1016] = -16'd256;
assign W_R_STAGE_LUT[1017] = 16'd3;
assign W_I_STAGE_LUT[1017] = -16'd256;
assign W_R_STAGE_LUT[1018] = 16'd2;
assign W_I_STAGE_LUT[1018] = -16'd256;
assign W_R_STAGE_LUT[1019] = 16'd2;
assign W_I_STAGE_LUT[1019] = -16'd256;
assign W_R_STAGE_LUT[1020] = 16'd2;
assign W_I_STAGE_LUT[1020] = -16'd256;
assign W_R_STAGE_LUT[1021] = 16'd1;
assign W_I_STAGE_LUT[1021] = -16'd256;
assign W_R_STAGE_LUT[1022] = 16'd1;
assign W_I_STAGE_LUT[1022] = -16'd256;
assign W_R_STAGE_LUT[1023] = 16'd0;
assign W_I_STAGE_LUT[1023] = -16'd256;
assign W_R_STAGE_LUT[1024] = 16'd0;
assign W_I_STAGE_LUT[1024] = -16'd256;
assign W_R_STAGE_LUT[1025] = 16'd0;
assign W_I_STAGE_LUT[1025] = -16'd256;
assign W_R_STAGE_LUT[1026] = -16'd1;
assign W_I_STAGE_LUT[1026] = -16'd256;
assign W_R_STAGE_LUT[1027] = -16'd1;
assign W_I_STAGE_LUT[1027] = -16'd256;
assign W_R_STAGE_LUT[1028] = -16'd2;
assign W_I_STAGE_LUT[1028] = -16'd256;
assign W_R_STAGE_LUT[1029] = -16'd2;
assign W_I_STAGE_LUT[1029] = -16'd256;
assign W_R_STAGE_LUT[1030] = -16'd2;
assign W_I_STAGE_LUT[1030] = -16'd256;
assign W_R_STAGE_LUT[1031] = -16'd3;
assign W_I_STAGE_LUT[1031] = -16'd256;
assign W_R_STAGE_LUT[1032] = -16'd3;
assign W_I_STAGE_LUT[1032] = -16'd256;
assign W_R_STAGE_LUT[1033] = -16'd4;
assign W_I_STAGE_LUT[1033] = -16'd256;
assign W_R_STAGE_LUT[1034] = -16'd4;
assign W_I_STAGE_LUT[1034] = -16'd256;
assign W_R_STAGE_LUT[1035] = -16'd4;
assign W_I_STAGE_LUT[1035] = -16'd256;
assign W_R_STAGE_LUT[1036] = -16'd5;
assign W_I_STAGE_LUT[1036] = -16'd256;
assign W_R_STAGE_LUT[1037] = -16'd5;
assign W_I_STAGE_LUT[1037] = -16'd256;
assign W_R_STAGE_LUT[1038] = -16'd5;
assign W_I_STAGE_LUT[1038] = -16'd256;
assign W_R_STAGE_LUT[1039] = -16'd6;
assign W_I_STAGE_LUT[1039] = -16'd256;
assign W_R_STAGE_LUT[1040] = -16'd6;
assign W_I_STAGE_LUT[1040] = -16'd256;
assign W_R_STAGE_LUT[1041] = -16'd7;
assign W_I_STAGE_LUT[1041] = -16'd256;
assign W_R_STAGE_LUT[1042] = -16'd7;
assign W_I_STAGE_LUT[1042] = -16'd256;
assign W_R_STAGE_LUT[1043] = -16'd7;
assign W_I_STAGE_LUT[1043] = -16'd256;
assign W_R_STAGE_LUT[1044] = -16'd8;
assign W_I_STAGE_LUT[1044] = -16'd256;
assign W_R_STAGE_LUT[1045] = -16'd8;
assign W_I_STAGE_LUT[1045] = -16'd256;
assign W_R_STAGE_LUT[1046] = -16'd9;
assign W_I_STAGE_LUT[1046] = -16'd256;
assign W_R_STAGE_LUT[1047] = -16'd9;
assign W_I_STAGE_LUT[1047] = -16'd256;
assign W_R_STAGE_LUT[1048] = -16'd9;
assign W_I_STAGE_LUT[1048] = -16'd256;
assign W_R_STAGE_LUT[1049] = -16'd10;
assign W_I_STAGE_LUT[1049] = -16'd256;
assign W_R_STAGE_LUT[1050] = -16'd10;
assign W_I_STAGE_LUT[1050] = -16'd256;
assign W_R_STAGE_LUT[1051] = -16'd11;
assign W_I_STAGE_LUT[1051] = -16'd256;
assign W_R_STAGE_LUT[1052] = -16'd11;
assign W_I_STAGE_LUT[1052] = -16'd256;
assign W_R_STAGE_LUT[1053] = -16'd11;
assign W_I_STAGE_LUT[1053] = -16'd256;
assign W_R_STAGE_LUT[1054] = -16'd12;
assign W_I_STAGE_LUT[1054] = -16'd256;
assign W_R_STAGE_LUT[1055] = -16'd12;
assign W_I_STAGE_LUT[1055] = -16'd256;
assign W_R_STAGE_LUT[1056] = -16'd13;
assign W_I_STAGE_LUT[1056] = -16'd256;
assign W_R_STAGE_LUT[1057] = -16'd13;
assign W_I_STAGE_LUT[1057] = -16'd256;
assign W_R_STAGE_LUT[1058] = -16'd13;
assign W_I_STAGE_LUT[1058] = -16'd256;
assign W_R_STAGE_LUT[1059] = -16'd14;
assign W_I_STAGE_LUT[1059] = -16'd256;
assign W_R_STAGE_LUT[1060] = -16'd14;
assign W_I_STAGE_LUT[1060] = -16'd256;
assign W_R_STAGE_LUT[1061] = -16'd15;
assign W_I_STAGE_LUT[1061] = -16'd256;
assign W_R_STAGE_LUT[1062] = -16'd15;
assign W_I_STAGE_LUT[1062] = -16'd256;
assign W_R_STAGE_LUT[1063] = -16'd15;
assign W_I_STAGE_LUT[1063] = -16'd256;
assign W_R_STAGE_LUT[1064] = -16'd16;
assign W_I_STAGE_LUT[1064] = -16'd256;
assign W_R_STAGE_LUT[1065] = -16'd16;
assign W_I_STAGE_LUT[1065] = -16'd255;
assign W_R_STAGE_LUT[1066] = -16'd16;
assign W_I_STAGE_LUT[1066] = -16'd255;
assign W_R_STAGE_LUT[1067] = -16'd17;
assign W_I_STAGE_LUT[1067] = -16'd255;
assign W_R_STAGE_LUT[1068] = -16'd17;
assign W_I_STAGE_LUT[1068] = -16'd255;
assign W_R_STAGE_LUT[1069] = -16'd18;
assign W_I_STAGE_LUT[1069] = -16'd255;
assign W_R_STAGE_LUT[1070] = -16'd18;
assign W_I_STAGE_LUT[1070] = -16'd255;
assign W_R_STAGE_LUT[1071] = -16'd18;
assign W_I_STAGE_LUT[1071] = -16'd255;
assign W_R_STAGE_LUT[1072] = -16'd19;
assign W_I_STAGE_LUT[1072] = -16'd255;
assign W_R_STAGE_LUT[1073] = -16'd19;
assign W_I_STAGE_LUT[1073] = -16'd255;
assign W_R_STAGE_LUT[1074] = -16'd20;
assign W_I_STAGE_LUT[1074] = -16'd255;
assign W_R_STAGE_LUT[1075] = -16'd20;
assign W_I_STAGE_LUT[1075] = -16'd255;
assign W_R_STAGE_LUT[1076] = -16'd20;
assign W_I_STAGE_LUT[1076] = -16'd255;
assign W_R_STAGE_LUT[1077] = -16'd21;
assign W_I_STAGE_LUT[1077] = -16'd255;
assign W_R_STAGE_LUT[1078] = -16'd21;
assign W_I_STAGE_LUT[1078] = -16'd255;
assign W_R_STAGE_LUT[1079] = -16'd22;
assign W_I_STAGE_LUT[1079] = -16'd255;
assign W_R_STAGE_LUT[1080] = -16'd22;
assign W_I_STAGE_LUT[1080] = -16'd255;
assign W_R_STAGE_LUT[1081] = -16'd22;
assign W_I_STAGE_LUT[1081] = -16'd255;
assign W_R_STAGE_LUT[1082] = -16'd23;
assign W_I_STAGE_LUT[1082] = -16'd255;
assign W_R_STAGE_LUT[1083] = -16'd23;
assign W_I_STAGE_LUT[1083] = -16'd255;
assign W_R_STAGE_LUT[1084] = -16'd24;
assign W_I_STAGE_LUT[1084] = -16'd255;
assign W_R_STAGE_LUT[1085] = -16'd24;
assign W_I_STAGE_LUT[1085] = -16'd255;
assign W_R_STAGE_LUT[1086] = -16'd24;
assign W_I_STAGE_LUT[1086] = -16'd255;
assign W_R_STAGE_LUT[1087] = -16'd25;
assign W_I_STAGE_LUT[1087] = -16'd255;
assign W_R_STAGE_LUT[1088] = -16'd25;
assign W_I_STAGE_LUT[1088] = -16'd255;
assign W_R_STAGE_LUT[1089] = -16'd25;
assign W_I_STAGE_LUT[1089] = -16'd255;
assign W_R_STAGE_LUT[1090] = -16'd26;
assign W_I_STAGE_LUT[1090] = -16'd255;
assign W_R_STAGE_LUT[1091] = -16'd26;
assign W_I_STAGE_LUT[1091] = -16'd255;
assign W_R_STAGE_LUT[1092] = -16'd27;
assign W_I_STAGE_LUT[1092] = -16'd255;
assign W_R_STAGE_LUT[1093] = -16'd27;
assign W_I_STAGE_LUT[1093] = -16'd255;
assign W_R_STAGE_LUT[1094] = -16'd27;
assign W_I_STAGE_LUT[1094] = -16'd255;
assign W_R_STAGE_LUT[1095] = -16'd28;
assign W_I_STAGE_LUT[1095] = -16'd254;
assign W_R_STAGE_LUT[1096] = -16'd28;
assign W_I_STAGE_LUT[1096] = -16'd254;
assign W_R_STAGE_LUT[1097] = -16'd29;
assign W_I_STAGE_LUT[1097] = -16'd254;
assign W_R_STAGE_LUT[1098] = -16'd29;
assign W_I_STAGE_LUT[1098] = -16'd254;
assign W_R_STAGE_LUT[1099] = -16'd29;
assign W_I_STAGE_LUT[1099] = -16'd254;
assign W_R_STAGE_LUT[1100] = -16'd30;
assign W_I_STAGE_LUT[1100] = -16'd254;
assign W_R_STAGE_LUT[1101] = -16'd30;
assign W_I_STAGE_LUT[1101] = -16'd254;
assign W_R_STAGE_LUT[1102] = -16'd31;
assign W_I_STAGE_LUT[1102] = -16'd254;
assign W_R_STAGE_LUT[1103] = -16'd31;
assign W_I_STAGE_LUT[1103] = -16'd254;
assign W_R_STAGE_LUT[1104] = -16'd31;
assign W_I_STAGE_LUT[1104] = -16'd254;
assign W_R_STAGE_LUT[1105] = -16'd32;
assign W_I_STAGE_LUT[1105] = -16'd254;
assign W_R_STAGE_LUT[1106] = -16'd32;
assign W_I_STAGE_LUT[1106] = -16'd254;
assign W_R_STAGE_LUT[1107] = -16'd33;
assign W_I_STAGE_LUT[1107] = -16'd254;
assign W_R_STAGE_LUT[1108] = -16'd33;
assign W_I_STAGE_LUT[1108] = -16'd254;
assign W_R_STAGE_LUT[1109] = -16'd33;
assign W_I_STAGE_LUT[1109] = -16'd254;
assign W_R_STAGE_LUT[1110] = -16'd34;
assign W_I_STAGE_LUT[1110] = -16'd254;
assign W_R_STAGE_LUT[1111] = -16'd34;
assign W_I_STAGE_LUT[1111] = -16'd254;
assign W_R_STAGE_LUT[1112] = -16'd34;
assign W_I_STAGE_LUT[1112] = -16'd254;
assign W_R_STAGE_LUT[1113] = -16'd35;
assign W_I_STAGE_LUT[1113] = -16'd254;
assign W_R_STAGE_LUT[1114] = -16'd35;
assign W_I_STAGE_LUT[1114] = -16'd254;
assign W_R_STAGE_LUT[1115] = -16'd36;
assign W_I_STAGE_LUT[1115] = -16'd254;
assign W_R_STAGE_LUT[1116] = -16'd36;
assign W_I_STAGE_LUT[1116] = -16'd253;
assign W_R_STAGE_LUT[1117] = -16'd36;
assign W_I_STAGE_LUT[1117] = -16'd253;
assign W_R_STAGE_LUT[1118] = -16'd37;
assign W_I_STAGE_LUT[1118] = -16'd253;
assign W_R_STAGE_LUT[1119] = -16'd37;
assign W_I_STAGE_LUT[1119] = -16'd253;
assign W_R_STAGE_LUT[1120] = -16'd38;
assign W_I_STAGE_LUT[1120] = -16'd253;
assign W_R_STAGE_LUT[1121] = -16'd38;
assign W_I_STAGE_LUT[1121] = -16'd253;
assign W_R_STAGE_LUT[1122] = -16'd38;
assign W_I_STAGE_LUT[1122] = -16'd253;
assign W_R_STAGE_LUT[1123] = -16'd39;
assign W_I_STAGE_LUT[1123] = -16'd253;
assign W_R_STAGE_LUT[1124] = -16'd39;
assign W_I_STAGE_LUT[1124] = -16'd253;
assign W_R_STAGE_LUT[1125] = -16'd40;
assign W_I_STAGE_LUT[1125] = -16'd253;
assign W_R_STAGE_LUT[1126] = -16'd40;
assign W_I_STAGE_LUT[1126] = -16'd253;
assign W_R_STAGE_LUT[1127] = -16'd40;
assign W_I_STAGE_LUT[1127] = -16'd253;
assign W_R_STAGE_LUT[1128] = -16'd41;
assign W_I_STAGE_LUT[1128] = -16'd253;
assign W_R_STAGE_LUT[1129] = -16'd41;
assign W_I_STAGE_LUT[1129] = -16'd253;
assign W_R_STAGE_LUT[1130] = -16'd41;
assign W_I_STAGE_LUT[1130] = -16'd253;
assign W_R_STAGE_LUT[1131] = -16'd42;
assign W_I_STAGE_LUT[1131] = -16'd253;
assign W_R_STAGE_LUT[1132] = -16'd42;
assign W_I_STAGE_LUT[1132] = -16'd252;
assign W_R_STAGE_LUT[1133] = -16'd43;
assign W_I_STAGE_LUT[1133] = -16'd252;
assign W_R_STAGE_LUT[1134] = -16'd43;
assign W_I_STAGE_LUT[1134] = -16'd252;
assign W_R_STAGE_LUT[1135] = -16'd43;
assign W_I_STAGE_LUT[1135] = -16'd252;
assign W_R_STAGE_LUT[1136] = -16'd44;
assign W_I_STAGE_LUT[1136] = -16'd252;
assign W_R_STAGE_LUT[1137] = -16'd44;
assign W_I_STAGE_LUT[1137] = -16'd252;
assign W_R_STAGE_LUT[1138] = -16'd45;
assign W_I_STAGE_LUT[1138] = -16'd252;
assign W_R_STAGE_LUT[1139] = -16'd45;
assign W_I_STAGE_LUT[1139] = -16'd252;
assign W_R_STAGE_LUT[1140] = -16'd45;
assign W_I_STAGE_LUT[1140] = -16'd252;
assign W_R_STAGE_LUT[1141] = -16'd46;
assign W_I_STAGE_LUT[1141] = -16'd252;
assign W_R_STAGE_LUT[1142] = -16'd46;
assign W_I_STAGE_LUT[1142] = -16'd252;
assign W_R_STAGE_LUT[1143] = -16'd46;
assign W_I_STAGE_LUT[1143] = -16'd252;
assign W_R_STAGE_LUT[1144] = -16'd47;
assign W_I_STAGE_LUT[1144] = -16'd252;
assign W_R_STAGE_LUT[1145] = -16'd47;
assign W_I_STAGE_LUT[1145] = -16'd252;
assign W_R_STAGE_LUT[1146] = -16'd48;
assign W_I_STAGE_LUT[1146] = -16'd252;
assign W_R_STAGE_LUT[1147] = -16'd48;
assign W_I_STAGE_LUT[1147] = -16'd251;
assign W_R_STAGE_LUT[1148] = -16'd48;
assign W_I_STAGE_LUT[1148] = -16'd251;
assign W_R_STAGE_LUT[1149] = -16'd49;
assign W_I_STAGE_LUT[1149] = -16'd251;
assign W_R_STAGE_LUT[1150] = -16'd49;
assign W_I_STAGE_LUT[1150] = -16'd251;
assign W_R_STAGE_LUT[1151] = -16'd50;
assign W_I_STAGE_LUT[1151] = -16'd251;
assign W_R_STAGE_LUT[1152] = -16'd50;
assign W_I_STAGE_LUT[1152] = -16'd251;
assign W_R_STAGE_LUT[1153] = -16'd50;
assign W_I_STAGE_LUT[1153] = -16'd251;
assign W_R_STAGE_LUT[1154] = -16'd51;
assign W_I_STAGE_LUT[1154] = -16'd251;
assign W_R_STAGE_LUT[1155] = -16'd51;
assign W_I_STAGE_LUT[1155] = -16'd251;
assign W_R_STAGE_LUT[1156] = -16'd51;
assign W_I_STAGE_LUT[1156] = -16'd251;
assign W_R_STAGE_LUT[1157] = -16'd52;
assign W_I_STAGE_LUT[1157] = -16'd251;
assign W_R_STAGE_LUT[1158] = -16'd52;
assign W_I_STAGE_LUT[1158] = -16'd251;
assign W_R_STAGE_LUT[1159] = -16'd53;
assign W_I_STAGE_LUT[1159] = -16'd251;
assign W_R_STAGE_LUT[1160] = -16'd53;
assign W_I_STAGE_LUT[1160] = -16'd250;
assign W_R_STAGE_LUT[1161] = -16'd53;
assign W_I_STAGE_LUT[1161] = -16'd250;
assign W_R_STAGE_LUT[1162] = -16'd54;
assign W_I_STAGE_LUT[1162] = -16'd250;
assign W_R_STAGE_LUT[1163] = -16'd54;
assign W_I_STAGE_LUT[1163] = -16'd250;
assign W_R_STAGE_LUT[1164] = -16'd55;
assign W_I_STAGE_LUT[1164] = -16'd250;
assign W_R_STAGE_LUT[1165] = -16'd55;
assign W_I_STAGE_LUT[1165] = -16'd250;
assign W_R_STAGE_LUT[1166] = -16'd55;
assign W_I_STAGE_LUT[1166] = -16'd250;
assign W_R_STAGE_LUT[1167] = -16'd56;
assign W_I_STAGE_LUT[1167] = -16'd250;
assign W_R_STAGE_LUT[1168] = -16'd56;
assign W_I_STAGE_LUT[1168] = -16'd250;
assign W_R_STAGE_LUT[1169] = -16'd56;
assign W_I_STAGE_LUT[1169] = -16'd250;
assign W_R_STAGE_LUT[1170] = -16'd57;
assign W_I_STAGE_LUT[1170] = -16'd250;
assign W_R_STAGE_LUT[1171] = -16'd57;
assign W_I_STAGE_LUT[1171] = -16'd250;
assign W_R_STAGE_LUT[1172] = -16'd58;
assign W_I_STAGE_LUT[1172] = -16'd249;
assign W_R_STAGE_LUT[1173] = -16'd58;
assign W_I_STAGE_LUT[1173] = -16'd249;
assign W_R_STAGE_LUT[1174] = -16'd58;
assign W_I_STAGE_LUT[1174] = -16'd249;
assign W_R_STAGE_LUT[1175] = -16'd59;
assign W_I_STAGE_LUT[1175] = -16'd249;
assign W_R_STAGE_LUT[1176] = -16'd59;
assign W_I_STAGE_LUT[1176] = -16'd249;
assign W_R_STAGE_LUT[1177] = -16'd60;
assign W_I_STAGE_LUT[1177] = -16'd249;
assign W_R_STAGE_LUT[1178] = -16'd60;
assign W_I_STAGE_LUT[1178] = -16'd249;
assign W_R_STAGE_LUT[1179] = -16'd60;
assign W_I_STAGE_LUT[1179] = -16'd249;
assign W_R_STAGE_LUT[1180] = -16'd61;
assign W_I_STAGE_LUT[1180] = -16'd249;
assign W_R_STAGE_LUT[1181] = -16'd61;
assign W_I_STAGE_LUT[1181] = -16'd249;
assign W_R_STAGE_LUT[1182] = -16'd61;
assign W_I_STAGE_LUT[1182] = -16'd249;
assign W_R_STAGE_LUT[1183] = -16'd62;
assign W_I_STAGE_LUT[1183] = -16'd248;
assign W_R_STAGE_LUT[1184] = -16'd62;
assign W_I_STAGE_LUT[1184] = -16'd248;
assign W_R_STAGE_LUT[1185] = -16'd63;
assign W_I_STAGE_LUT[1185] = -16'd248;
assign W_R_STAGE_LUT[1186] = -16'd63;
assign W_I_STAGE_LUT[1186] = -16'd248;
assign W_R_STAGE_LUT[1187] = -16'd63;
assign W_I_STAGE_LUT[1187] = -16'd248;
assign W_R_STAGE_LUT[1188] = -16'd64;
assign W_I_STAGE_LUT[1188] = -16'd248;
assign W_R_STAGE_LUT[1189] = -16'd64;
assign W_I_STAGE_LUT[1189] = -16'd248;
assign W_R_STAGE_LUT[1190] = -16'd64;
assign W_I_STAGE_LUT[1190] = -16'd248;
assign W_R_STAGE_LUT[1191] = -16'd65;
assign W_I_STAGE_LUT[1191] = -16'd248;
assign W_R_STAGE_LUT[1192] = -16'd65;
assign W_I_STAGE_LUT[1192] = -16'd248;
assign W_R_STAGE_LUT[1193] = -16'd66;
assign W_I_STAGE_LUT[1193] = -16'd247;
assign W_R_STAGE_LUT[1194] = -16'd66;
assign W_I_STAGE_LUT[1194] = -16'd247;
assign W_R_STAGE_LUT[1195] = -16'd66;
assign W_I_STAGE_LUT[1195] = -16'd247;
assign W_R_STAGE_LUT[1196] = -16'd67;
assign W_I_STAGE_LUT[1196] = -16'd247;
assign W_R_STAGE_LUT[1197] = -16'd67;
assign W_I_STAGE_LUT[1197] = -16'd247;
assign W_R_STAGE_LUT[1198] = -16'd68;
assign W_I_STAGE_LUT[1198] = -16'd247;
assign W_R_STAGE_LUT[1199] = -16'd68;
assign W_I_STAGE_LUT[1199] = -16'd247;
assign W_R_STAGE_LUT[1200] = -16'd68;
assign W_I_STAGE_LUT[1200] = -16'd247;
assign W_R_STAGE_LUT[1201] = -16'd69;
assign W_I_STAGE_LUT[1201] = -16'd247;
assign W_R_STAGE_LUT[1202] = -16'd69;
assign W_I_STAGE_LUT[1202] = -16'd247;
assign W_R_STAGE_LUT[1203] = -16'd69;
assign W_I_STAGE_LUT[1203] = -16'd246;
assign W_R_STAGE_LUT[1204] = -16'd70;
assign W_I_STAGE_LUT[1204] = -16'd246;
assign W_R_STAGE_LUT[1205] = -16'd70;
assign W_I_STAGE_LUT[1205] = -16'd246;
assign W_R_STAGE_LUT[1206] = -16'd71;
assign W_I_STAGE_LUT[1206] = -16'd246;
assign W_R_STAGE_LUT[1207] = -16'd71;
assign W_I_STAGE_LUT[1207] = -16'd246;
assign W_R_STAGE_LUT[1208] = -16'd71;
assign W_I_STAGE_LUT[1208] = -16'd246;
assign W_R_STAGE_LUT[1209] = -16'd72;
assign W_I_STAGE_LUT[1209] = -16'd246;
assign W_R_STAGE_LUT[1210] = -16'd72;
assign W_I_STAGE_LUT[1210] = -16'd246;
assign W_R_STAGE_LUT[1211] = -16'd72;
assign W_I_STAGE_LUT[1211] = -16'd246;
assign W_R_STAGE_LUT[1212] = -16'd73;
assign W_I_STAGE_LUT[1212] = -16'd245;
assign W_R_STAGE_LUT[1213] = -16'd73;
assign W_I_STAGE_LUT[1213] = -16'd245;
assign W_R_STAGE_LUT[1214] = -16'd74;
assign W_I_STAGE_LUT[1214] = -16'd245;
assign W_R_STAGE_LUT[1215] = -16'd74;
assign W_I_STAGE_LUT[1215] = -16'd245;
assign W_R_STAGE_LUT[1216] = -16'd74;
assign W_I_STAGE_LUT[1216] = -16'd245;
assign W_R_STAGE_LUT[1217] = -16'd75;
assign W_I_STAGE_LUT[1217] = -16'd245;
assign W_R_STAGE_LUT[1218] = -16'd75;
assign W_I_STAGE_LUT[1218] = -16'd245;
assign W_R_STAGE_LUT[1219] = -16'd75;
assign W_I_STAGE_LUT[1219] = -16'd245;
assign W_R_STAGE_LUT[1220] = -16'd76;
assign W_I_STAGE_LUT[1220] = -16'd245;
assign W_R_STAGE_LUT[1221] = -16'd76;
assign W_I_STAGE_LUT[1221] = -16'd244;
assign W_R_STAGE_LUT[1222] = -16'd77;
assign W_I_STAGE_LUT[1222] = -16'd244;
assign W_R_STAGE_LUT[1223] = -16'd77;
assign W_I_STAGE_LUT[1223] = -16'd244;
assign W_R_STAGE_LUT[1224] = -16'd77;
assign W_I_STAGE_LUT[1224] = -16'd244;
assign W_R_STAGE_LUT[1225] = -16'd78;
assign W_I_STAGE_LUT[1225] = -16'd244;
assign W_R_STAGE_LUT[1226] = -16'd78;
assign W_I_STAGE_LUT[1226] = -16'd244;
assign W_R_STAGE_LUT[1227] = -16'd78;
assign W_I_STAGE_LUT[1227] = -16'd244;
assign W_R_STAGE_LUT[1228] = -16'd79;
assign W_I_STAGE_LUT[1228] = -16'd244;
assign W_R_STAGE_LUT[1229] = -16'd79;
assign W_I_STAGE_LUT[1229] = -16'd243;
assign W_R_STAGE_LUT[1230] = -16'd80;
assign W_I_STAGE_LUT[1230] = -16'd243;
assign W_R_STAGE_LUT[1231] = -16'd80;
assign W_I_STAGE_LUT[1231] = -16'd243;
assign W_R_STAGE_LUT[1232] = -16'd80;
assign W_I_STAGE_LUT[1232] = -16'd243;
assign W_R_STAGE_LUT[1233] = -16'd81;
assign W_I_STAGE_LUT[1233] = -16'd243;
assign W_R_STAGE_LUT[1234] = -16'd81;
assign W_I_STAGE_LUT[1234] = -16'd243;
assign W_R_STAGE_LUT[1235] = -16'd81;
assign W_I_STAGE_LUT[1235] = -16'd243;
assign W_R_STAGE_LUT[1236] = -16'd82;
assign W_I_STAGE_LUT[1236] = -16'd243;
assign W_R_STAGE_LUT[1237] = -16'd82;
assign W_I_STAGE_LUT[1237] = -16'd242;
assign W_R_STAGE_LUT[1238] = -16'd83;
assign W_I_STAGE_LUT[1238] = -16'd242;
assign W_R_STAGE_LUT[1239] = -16'd83;
assign W_I_STAGE_LUT[1239] = -16'd242;
assign W_R_STAGE_LUT[1240] = -16'd83;
assign W_I_STAGE_LUT[1240] = -16'd242;
assign W_R_STAGE_LUT[1241] = -16'd84;
assign W_I_STAGE_LUT[1241] = -16'd242;
assign W_R_STAGE_LUT[1242] = -16'd84;
assign W_I_STAGE_LUT[1242] = -16'd242;
assign W_R_STAGE_LUT[1243] = -16'd84;
assign W_I_STAGE_LUT[1243] = -16'd242;
assign W_R_STAGE_LUT[1244] = -16'd85;
assign W_I_STAGE_LUT[1244] = -16'd242;
assign W_R_STAGE_LUT[1245] = -16'd85;
assign W_I_STAGE_LUT[1245] = -16'd241;
assign W_R_STAGE_LUT[1246] = -16'd86;
assign W_I_STAGE_LUT[1246] = -16'd241;
assign W_R_STAGE_LUT[1247] = -16'd86;
assign W_I_STAGE_LUT[1247] = -16'd241;
assign W_R_STAGE_LUT[1248] = -16'd86;
assign W_I_STAGE_LUT[1248] = -16'd241;
assign W_R_STAGE_LUT[1249] = -16'd87;
assign W_I_STAGE_LUT[1249] = -16'd241;
assign W_R_STAGE_LUT[1250] = -16'd87;
assign W_I_STAGE_LUT[1250] = -16'd241;
assign W_R_STAGE_LUT[1251] = -16'd87;
assign W_I_STAGE_LUT[1251] = -16'd241;
assign W_R_STAGE_LUT[1252] = -16'd88;
assign W_I_STAGE_LUT[1252] = -16'd241;
assign W_R_STAGE_LUT[1253] = -16'd88;
assign W_I_STAGE_LUT[1253] = -16'd240;
assign W_R_STAGE_LUT[1254] = -16'd88;
assign W_I_STAGE_LUT[1254] = -16'd240;
assign W_R_STAGE_LUT[1255] = -16'd89;
assign W_I_STAGE_LUT[1255] = -16'd240;
assign W_R_STAGE_LUT[1256] = -16'd89;
assign W_I_STAGE_LUT[1256] = -16'd240;
assign W_R_STAGE_LUT[1257] = -16'd90;
assign W_I_STAGE_LUT[1257] = -16'd240;
assign W_R_STAGE_LUT[1258] = -16'd90;
assign W_I_STAGE_LUT[1258] = -16'd240;
assign W_R_STAGE_LUT[1259] = -16'd90;
assign W_I_STAGE_LUT[1259] = -16'd240;
assign W_R_STAGE_LUT[1260] = -16'd91;
assign W_I_STAGE_LUT[1260] = -16'd239;
assign W_R_STAGE_LUT[1261] = -16'd91;
assign W_I_STAGE_LUT[1261] = -16'd239;
assign W_R_STAGE_LUT[1262] = -16'd91;
assign W_I_STAGE_LUT[1262] = -16'd239;
assign W_R_STAGE_LUT[1263] = -16'd92;
assign W_I_STAGE_LUT[1263] = -16'd239;
assign W_R_STAGE_LUT[1264] = -16'd92;
assign W_I_STAGE_LUT[1264] = -16'd239;
assign W_R_STAGE_LUT[1265] = -16'd92;
assign W_I_STAGE_LUT[1265] = -16'd239;
assign W_R_STAGE_LUT[1266] = -16'd93;
assign W_I_STAGE_LUT[1266] = -16'd239;
assign W_R_STAGE_LUT[1267] = -16'd93;
assign W_I_STAGE_LUT[1267] = -16'd238;
assign W_R_STAGE_LUT[1268] = -16'd94;
assign W_I_STAGE_LUT[1268] = -16'd238;
assign W_R_STAGE_LUT[1269] = -16'd94;
assign W_I_STAGE_LUT[1269] = -16'd238;
assign W_R_STAGE_LUT[1270] = -16'd94;
assign W_I_STAGE_LUT[1270] = -16'd238;
assign W_R_STAGE_LUT[1271] = -16'd95;
assign W_I_STAGE_LUT[1271] = -16'd238;
assign W_R_STAGE_LUT[1272] = -16'd95;
assign W_I_STAGE_LUT[1272] = -16'd238;
assign W_R_STAGE_LUT[1273] = -16'd95;
assign W_I_STAGE_LUT[1273] = -16'd238;
assign W_R_STAGE_LUT[1274] = -16'd96;
assign W_I_STAGE_LUT[1274] = -16'd237;
assign W_R_STAGE_LUT[1275] = -16'd96;
assign W_I_STAGE_LUT[1275] = -16'd237;
assign W_R_STAGE_LUT[1276] = -16'd97;
assign W_I_STAGE_LUT[1276] = -16'd237;
assign W_R_STAGE_LUT[1277] = -16'd97;
assign W_I_STAGE_LUT[1277] = -16'd237;
assign W_R_STAGE_LUT[1278] = -16'd97;
assign W_I_STAGE_LUT[1278] = -16'd237;
assign W_R_STAGE_LUT[1279] = -16'd98;
assign W_I_STAGE_LUT[1279] = -16'd237;
assign W_R_STAGE_LUT[1280] = -16'd98;
assign W_I_STAGE_LUT[1280] = -16'd237;
assign W_R_STAGE_LUT[1281] = -16'd98;
assign W_I_STAGE_LUT[1281] = -16'd236;
assign W_R_STAGE_LUT[1282] = -16'd99;
assign W_I_STAGE_LUT[1282] = -16'd236;
assign W_R_STAGE_LUT[1283] = -16'd99;
assign W_I_STAGE_LUT[1283] = -16'd236;
assign W_R_STAGE_LUT[1284] = -16'd99;
assign W_I_STAGE_LUT[1284] = -16'd236;
assign W_R_STAGE_LUT[1285] = -16'd100;
assign W_I_STAGE_LUT[1285] = -16'd236;
assign W_R_STAGE_LUT[1286] = -16'd100;
assign W_I_STAGE_LUT[1286] = -16'd236;
assign W_R_STAGE_LUT[1287] = -16'd101;
assign W_I_STAGE_LUT[1287] = -16'd235;
assign W_R_STAGE_LUT[1288] = -16'd101;
assign W_I_STAGE_LUT[1288] = -16'd235;
assign W_R_STAGE_LUT[1289] = -16'd101;
assign W_I_STAGE_LUT[1289] = -16'd235;
assign W_R_STAGE_LUT[1290] = -16'd102;
assign W_I_STAGE_LUT[1290] = -16'd235;
assign W_R_STAGE_LUT[1291] = -16'd102;
assign W_I_STAGE_LUT[1291] = -16'd235;
assign W_R_STAGE_LUT[1292] = -16'd102;
assign W_I_STAGE_LUT[1292] = -16'd235;
assign W_R_STAGE_LUT[1293] = -16'd103;
assign W_I_STAGE_LUT[1293] = -16'd235;
assign W_R_STAGE_LUT[1294] = -16'd103;
assign W_I_STAGE_LUT[1294] = -16'd234;
assign W_R_STAGE_LUT[1295] = -16'd103;
assign W_I_STAGE_LUT[1295] = -16'd234;
assign W_R_STAGE_LUT[1296] = -16'd104;
assign W_I_STAGE_LUT[1296] = -16'd234;
assign W_R_STAGE_LUT[1297] = -16'd104;
assign W_I_STAGE_LUT[1297] = -16'd234;
assign W_R_STAGE_LUT[1298] = -16'd104;
assign W_I_STAGE_LUT[1298] = -16'd234;
assign W_R_STAGE_LUT[1299] = -16'd105;
assign W_I_STAGE_LUT[1299] = -16'd234;
assign W_R_STAGE_LUT[1300] = -16'd105;
assign W_I_STAGE_LUT[1300] = -16'd233;
assign W_R_STAGE_LUT[1301] = -16'd106;
assign W_I_STAGE_LUT[1301] = -16'd233;
assign W_R_STAGE_LUT[1302] = -16'd106;
assign W_I_STAGE_LUT[1302] = -16'd233;
assign W_R_STAGE_LUT[1303] = -16'd106;
assign W_I_STAGE_LUT[1303] = -16'd233;
assign W_R_STAGE_LUT[1304] = -16'd107;
assign W_I_STAGE_LUT[1304] = -16'd233;
assign W_R_STAGE_LUT[1305] = -16'd107;
assign W_I_STAGE_LUT[1305] = -16'd233;
assign W_R_STAGE_LUT[1306] = -16'd107;
assign W_I_STAGE_LUT[1306] = -16'd232;
assign W_R_STAGE_LUT[1307] = -16'd108;
assign W_I_STAGE_LUT[1307] = -16'd232;
assign W_R_STAGE_LUT[1308] = -16'd108;
assign W_I_STAGE_LUT[1308] = -16'd232;
assign W_R_STAGE_LUT[1309] = -16'd108;
assign W_I_STAGE_LUT[1309] = -16'd232;
assign W_R_STAGE_LUT[1310] = -16'd109;
assign W_I_STAGE_LUT[1310] = -16'd232;
assign W_R_STAGE_LUT[1311] = -16'd109;
assign W_I_STAGE_LUT[1311] = -16'd232;
assign W_R_STAGE_LUT[1312] = -16'd109;
assign W_I_STAGE_LUT[1312] = -16'd231;
assign W_R_STAGE_LUT[1313] = -16'd110;
assign W_I_STAGE_LUT[1313] = -16'd231;
assign W_R_STAGE_LUT[1314] = -16'd110;
assign W_I_STAGE_LUT[1314] = -16'd231;
assign W_R_STAGE_LUT[1315] = -16'd111;
assign W_I_STAGE_LUT[1315] = -16'd231;
assign W_R_STAGE_LUT[1316] = -16'd111;
assign W_I_STAGE_LUT[1316] = -16'd231;
assign W_R_STAGE_LUT[1317] = -16'd111;
assign W_I_STAGE_LUT[1317] = -16'd231;
assign W_R_STAGE_LUT[1318] = -16'd112;
assign W_I_STAGE_LUT[1318] = -16'd230;
assign W_R_STAGE_LUT[1319] = -16'd112;
assign W_I_STAGE_LUT[1319] = -16'd230;
assign W_R_STAGE_LUT[1320] = -16'd112;
assign W_I_STAGE_LUT[1320] = -16'd230;
assign W_R_STAGE_LUT[1321] = -16'd113;
assign W_I_STAGE_LUT[1321] = -16'd230;
assign W_R_STAGE_LUT[1322] = -16'd113;
assign W_I_STAGE_LUT[1322] = -16'd230;
assign W_R_STAGE_LUT[1323] = -16'd113;
assign W_I_STAGE_LUT[1323] = -16'd230;
assign W_R_STAGE_LUT[1324] = -16'd114;
assign W_I_STAGE_LUT[1324] = -16'd229;
assign W_R_STAGE_LUT[1325] = -16'd114;
assign W_I_STAGE_LUT[1325] = -16'd229;
assign W_R_STAGE_LUT[1326] = -16'd114;
assign W_I_STAGE_LUT[1326] = -16'd229;
assign W_R_STAGE_LUT[1327] = -16'd115;
assign W_I_STAGE_LUT[1327] = -16'd229;
assign W_R_STAGE_LUT[1328] = -16'd115;
assign W_I_STAGE_LUT[1328] = -16'd229;
assign W_R_STAGE_LUT[1329] = -16'd115;
assign W_I_STAGE_LUT[1329] = -16'd228;
assign W_R_STAGE_LUT[1330] = -16'd116;
assign W_I_STAGE_LUT[1330] = -16'd228;
assign W_R_STAGE_LUT[1331] = -16'd116;
assign W_I_STAGE_LUT[1331] = -16'd228;
assign W_R_STAGE_LUT[1332] = -16'd117;
assign W_I_STAGE_LUT[1332] = -16'd228;
assign W_R_STAGE_LUT[1333] = -16'd117;
assign W_I_STAGE_LUT[1333] = -16'd228;
assign W_R_STAGE_LUT[1334] = -16'd117;
assign W_I_STAGE_LUT[1334] = -16'd228;
assign W_R_STAGE_LUT[1335] = -16'd118;
assign W_I_STAGE_LUT[1335] = -16'd227;
assign W_R_STAGE_LUT[1336] = -16'd118;
assign W_I_STAGE_LUT[1336] = -16'd227;
assign W_R_STAGE_LUT[1337] = -16'd118;
assign W_I_STAGE_LUT[1337] = -16'd227;
assign W_R_STAGE_LUT[1338] = -16'd119;
assign W_I_STAGE_LUT[1338] = -16'd227;
assign W_R_STAGE_LUT[1339] = -16'd119;
assign W_I_STAGE_LUT[1339] = -16'd227;
assign W_R_STAGE_LUT[1340] = -16'd119;
assign W_I_STAGE_LUT[1340] = -16'd227;
assign W_R_STAGE_LUT[1341] = -16'd120;
assign W_I_STAGE_LUT[1341] = -16'd226;
assign W_R_STAGE_LUT[1342] = -16'd120;
assign W_I_STAGE_LUT[1342] = -16'd226;
assign W_R_STAGE_LUT[1343] = -16'd120;
assign W_I_STAGE_LUT[1343] = -16'd226;
assign W_R_STAGE_LUT[1344] = -16'd121;
assign W_I_STAGE_LUT[1344] = -16'd226;
assign W_R_STAGE_LUT[1345] = -16'd121;
assign W_I_STAGE_LUT[1345] = -16'd226;
assign W_R_STAGE_LUT[1346] = -16'd121;
assign W_I_STAGE_LUT[1346] = -16'd225;
assign W_R_STAGE_LUT[1347] = -16'd122;
assign W_I_STAGE_LUT[1347] = -16'd225;
assign W_R_STAGE_LUT[1348] = -16'd122;
assign W_I_STAGE_LUT[1348] = -16'd225;
assign W_R_STAGE_LUT[1349] = -16'd122;
assign W_I_STAGE_LUT[1349] = -16'd225;
assign W_R_STAGE_LUT[1350] = -16'd123;
assign W_I_STAGE_LUT[1350] = -16'd225;
assign W_R_STAGE_LUT[1351] = -16'd123;
assign W_I_STAGE_LUT[1351] = -16'd224;
assign W_R_STAGE_LUT[1352] = -16'd123;
assign W_I_STAGE_LUT[1352] = -16'd224;
assign W_R_STAGE_LUT[1353] = -16'd124;
assign W_I_STAGE_LUT[1353] = -16'd224;
assign W_R_STAGE_LUT[1354] = -16'd124;
assign W_I_STAGE_LUT[1354] = -16'd224;
assign W_R_STAGE_LUT[1355] = -16'd124;
assign W_I_STAGE_LUT[1355] = -16'd224;
assign W_R_STAGE_LUT[1356] = -16'd125;
assign W_I_STAGE_LUT[1356] = -16'd224;
assign W_R_STAGE_LUT[1357] = -16'd125;
assign W_I_STAGE_LUT[1357] = -16'd223;
assign W_R_STAGE_LUT[1358] = -16'd125;
assign W_I_STAGE_LUT[1358] = -16'd223;
assign W_R_STAGE_LUT[1359] = -16'd126;
assign W_I_STAGE_LUT[1359] = -16'd223;
assign W_R_STAGE_LUT[1360] = -16'd126;
assign W_I_STAGE_LUT[1360] = -16'd223;
assign W_R_STAGE_LUT[1361] = -16'd127;
assign W_I_STAGE_LUT[1361] = -16'd223;
assign W_R_STAGE_LUT[1362] = -16'd127;
assign W_I_STAGE_LUT[1362] = -16'd222;
assign W_R_STAGE_LUT[1363] = -16'd127;
assign W_I_STAGE_LUT[1363] = -16'd222;
assign W_R_STAGE_LUT[1364] = -16'd128;
assign W_I_STAGE_LUT[1364] = -16'd222;
assign W_R_STAGE_LUT[1365] = -16'd128;
assign W_I_STAGE_LUT[1365] = -16'd222;
assign W_R_STAGE_LUT[1366] = -16'd128;
assign W_I_STAGE_LUT[1366] = -16'd222;
assign W_R_STAGE_LUT[1367] = -16'd129;
assign W_I_STAGE_LUT[1367] = -16'd221;
assign W_R_STAGE_LUT[1368] = -16'd129;
assign W_I_STAGE_LUT[1368] = -16'd221;
assign W_R_STAGE_LUT[1369] = -16'd129;
assign W_I_STAGE_LUT[1369] = -16'd221;
assign W_R_STAGE_LUT[1370] = -16'd130;
assign W_I_STAGE_LUT[1370] = -16'd221;
assign W_R_STAGE_LUT[1371] = -16'd130;
assign W_I_STAGE_LUT[1371] = -16'd221;
assign W_R_STAGE_LUT[1372] = -16'd130;
assign W_I_STAGE_LUT[1372] = -16'd220;
assign W_R_STAGE_LUT[1373] = -16'd131;
assign W_I_STAGE_LUT[1373] = -16'd220;
assign W_R_STAGE_LUT[1374] = -16'd131;
assign W_I_STAGE_LUT[1374] = -16'd220;
assign W_R_STAGE_LUT[1375] = -16'd131;
assign W_I_STAGE_LUT[1375] = -16'd220;
assign W_R_STAGE_LUT[1376] = -16'd132;
assign W_I_STAGE_LUT[1376] = -16'd220;
assign W_R_STAGE_LUT[1377] = -16'd132;
assign W_I_STAGE_LUT[1377] = -16'd219;
assign W_R_STAGE_LUT[1378] = -16'd132;
assign W_I_STAGE_LUT[1378] = -16'd219;
assign W_R_STAGE_LUT[1379] = -16'd133;
assign W_I_STAGE_LUT[1379] = -16'd219;
assign W_R_STAGE_LUT[1380] = -16'd133;
assign W_I_STAGE_LUT[1380] = -16'd219;
assign W_R_STAGE_LUT[1381] = -16'd133;
assign W_I_STAGE_LUT[1381] = -16'd219;
assign W_R_STAGE_LUT[1382] = -16'd134;
assign W_I_STAGE_LUT[1382] = -16'd218;
assign W_R_STAGE_LUT[1383] = -16'd134;
assign W_I_STAGE_LUT[1383] = -16'd218;
assign W_R_STAGE_LUT[1384] = -16'd134;
assign W_I_STAGE_LUT[1384] = -16'd218;
assign W_R_STAGE_LUT[1385] = -16'd135;
assign W_I_STAGE_LUT[1385] = -16'd218;
assign W_R_STAGE_LUT[1386] = -16'd135;
assign W_I_STAGE_LUT[1386] = -16'd218;
assign W_R_STAGE_LUT[1387] = -16'd135;
assign W_I_STAGE_LUT[1387] = -16'd217;
assign W_R_STAGE_LUT[1388] = -16'd136;
assign W_I_STAGE_LUT[1388] = -16'd217;
assign W_R_STAGE_LUT[1389] = -16'd136;
assign W_I_STAGE_LUT[1389] = -16'd217;
assign W_R_STAGE_LUT[1390] = -16'd136;
assign W_I_STAGE_LUT[1390] = -16'd217;
assign W_R_STAGE_LUT[1391] = -16'd137;
assign W_I_STAGE_LUT[1391] = -16'd216;
assign W_R_STAGE_LUT[1392] = -16'd137;
assign W_I_STAGE_LUT[1392] = -16'd216;
assign W_R_STAGE_LUT[1393] = -16'd137;
assign W_I_STAGE_LUT[1393] = -16'd216;
assign W_R_STAGE_LUT[1394] = -16'd138;
assign W_I_STAGE_LUT[1394] = -16'd216;
assign W_R_STAGE_LUT[1395] = -16'd138;
assign W_I_STAGE_LUT[1395] = -16'd216;
assign W_R_STAGE_LUT[1396] = -16'd138;
assign W_I_STAGE_LUT[1396] = -16'd215;
assign W_R_STAGE_LUT[1397] = -16'd139;
assign W_I_STAGE_LUT[1397] = -16'd215;
assign W_R_STAGE_LUT[1398] = -16'd139;
assign W_I_STAGE_LUT[1398] = -16'd215;
assign W_R_STAGE_LUT[1399] = -16'd139;
assign W_I_STAGE_LUT[1399] = -16'd215;
assign W_R_STAGE_LUT[1400] = -16'd140;
assign W_I_STAGE_LUT[1400] = -16'd215;
assign W_R_STAGE_LUT[1401] = -16'd140;
assign W_I_STAGE_LUT[1401] = -16'd214;
assign W_R_STAGE_LUT[1402] = -16'd140;
assign W_I_STAGE_LUT[1402] = -16'd214;
assign W_R_STAGE_LUT[1403] = -16'd141;
assign W_I_STAGE_LUT[1403] = -16'd214;
assign W_R_STAGE_LUT[1404] = -16'd141;
assign W_I_STAGE_LUT[1404] = -16'd214;
assign W_R_STAGE_LUT[1405] = -16'd141;
assign W_I_STAGE_LUT[1405] = -16'd214;
assign W_R_STAGE_LUT[1406] = -16'd142;
assign W_I_STAGE_LUT[1406] = -16'd213;
assign W_R_STAGE_LUT[1407] = -16'd142;
assign W_I_STAGE_LUT[1407] = -16'd213;
assign W_R_STAGE_LUT[1408] = -16'd142;
assign W_I_STAGE_LUT[1408] = -16'd213;
assign W_R_STAGE_LUT[1409] = -16'd143;
assign W_I_STAGE_LUT[1409] = -16'd213;
assign W_R_STAGE_LUT[1410] = -16'd143;
assign W_I_STAGE_LUT[1410] = -16'd212;
assign W_R_STAGE_LUT[1411] = -16'd143;
assign W_I_STAGE_LUT[1411] = -16'd212;
assign W_R_STAGE_LUT[1412] = -16'd144;
assign W_I_STAGE_LUT[1412] = -16'd212;
assign W_R_STAGE_LUT[1413] = -16'd144;
assign W_I_STAGE_LUT[1413] = -16'd212;
assign W_R_STAGE_LUT[1414] = -16'd144;
assign W_I_STAGE_LUT[1414] = -16'd212;
assign W_R_STAGE_LUT[1415] = -16'd145;
assign W_I_STAGE_LUT[1415] = -16'd211;
assign W_R_STAGE_LUT[1416] = -16'd145;
assign W_I_STAGE_LUT[1416] = -16'd211;
assign W_R_STAGE_LUT[1417] = -16'd145;
assign W_I_STAGE_LUT[1417] = -16'd211;
assign W_R_STAGE_LUT[1418] = -16'd145;
assign W_I_STAGE_LUT[1418] = -16'd211;
assign W_R_STAGE_LUT[1419] = -16'd146;
assign W_I_STAGE_LUT[1419] = -16'd210;
assign W_R_STAGE_LUT[1420] = -16'd146;
assign W_I_STAGE_LUT[1420] = -16'd210;
assign W_R_STAGE_LUT[1421] = -16'd146;
assign W_I_STAGE_LUT[1421] = -16'd210;
assign W_R_STAGE_LUT[1422] = -16'd147;
assign W_I_STAGE_LUT[1422] = -16'd210;
assign W_R_STAGE_LUT[1423] = -16'd147;
assign W_I_STAGE_LUT[1423] = -16'd210;
assign W_R_STAGE_LUT[1424] = -16'd147;
assign W_I_STAGE_LUT[1424] = -16'd209;
assign W_R_STAGE_LUT[1425] = -16'd148;
assign W_I_STAGE_LUT[1425] = -16'd209;
assign W_R_STAGE_LUT[1426] = -16'd148;
assign W_I_STAGE_LUT[1426] = -16'd209;
assign W_R_STAGE_LUT[1427] = -16'd148;
assign W_I_STAGE_LUT[1427] = -16'd209;
assign W_R_STAGE_LUT[1428] = -16'd149;
assign W_I_STAGE_LUT[1428] = -16'd208;
assign W_R_STAGE_LUT[1429] = -16'd149;
assign W_I_STAGE_LUT[1429] = -16'd208;
assign W_R_STAGE_LUT[1430] = -16'd149;
assign W_I_STAGE_LUT[1430] = -16'd208;
assign W_R_STAGE_LUT[1431] = -16'd150;
assign W_I_STAGE_LUT[1431] = -16'd208;
assign W_R_STAGE_LUT[1432] = -16'd150;
assign W_I_STAGE_LUT[1432] = -16'd207;
assign W_R_STAGE_LUT[1433] = -16'd150;
assign W_I_STAGE_LUT[1433] = -16'd207;
assign W_R_STAGE_LUT[1434] = -16'd151;
assign W_I_STAGE_LUT[1434] = -16'd207;
assign W_R_STAGE_LUT[1435] = -16'd151;
assign W_I_STAGE_LUT[1435] = -16'd207;
assign W_R_STAGE_LUT[1436] = -16'd151;
assign W_I_STAGE_LUT[1436] = -16'd207;
assign W_R_STAGE_LUT[1437] = -16'd152;
assign W_I_STAGE_LUT[1437] = -16'd206;
assign W_R_STAGE_LUT[1438] = -16'd152;
assign W_I_STAGE_LUT[1438] = -16'd206;
assign W_R_STAGE_LUT[1439] = -16'd152;
assign W_I_STAGE_LUT[1439] = -16'd206;
assign W_R_STAGE_LUT[1440] = -16'd152;
assign W_I_STAGE_LUT[1440] = -16'd206;
assign W_R_STAGE_LUT[1441] = -16'd153;
assign W_I_STAGE_LUT[1441] = -16'd205;
assign W_R_STAGE_LUT[1442] = -16'd153;
assign W_I_STAGE_LUT[1442] = -16'd205;
assign W_R_STAGE_LUT[1443] = -16'd153;
assign W_I_STAGE_LUT[1443] = -16'd205;
assign W_R_STAGE_LUT[1444] = -16'd154;
assign W_I_STAGE_LUT[1444] = -16'd205;
assign W_R_STAGE_LUT[1445] = -16'd154;
assign W_I_STAGE_LUT[1445] = -16'd204;
assign W_R_STAGE_LUT[1446] = -16'd154;
assign W_I_STAGE_LUT[1446] = -16'd204;
assign W_R_STAGE_LUT[1447] = -16'd155;
assign W_I_STAGE_LUT[1447] = -16'd204;
assign W_R_STAGE_LUT[1448] = -16'd155;
assign W_I_STAGE_LUT[1448] = -16'd204;
assign W_R_STAGE_LUT[1449] = -16'd155;
assign W_I_STAGE_LUT[1449] = -16'd203;
assign W_R_STAGE_LUT[1450] = -16'd156;
assign W_I_STAGE_LUT[1450] = -16'd203;
assign W_R_STAGE_LUT[1451] = -16'd156;
assign W_I_STAGE_LUT[1451] = -16'd203;
assign W_R_STAGE_LUT[1452] = -16'd156;
assign W_I_STAGE_LUT[1452] = -16'd203;
assign W_R_STAGE_LUT[1453] = -16'd157;
assign W_I_STAGE_LUT[1453] = -16'd203;
assign W_R_STAGE_LUT[1454] = -16'd157;
assign W_I_STAGE_LUT[1454] = -16'd202;
assign W_R_STAGE_LUT[1455] = -16'd157;
assign W_I_STAGE_LUT[1455] = -16'd202;
assign W_R_STAGE_LUT[1456] = -16'd157;
assign W_I_STAGE_LUT[1456] = -16'd202;
assign W_R_STAGE_LUT[1457] = -16'd158;
assign W_I_STAGE_LUT[1457] = -16'd202;
assign W_R_STAGE_LUT[1458] = -16'd158;
assign W_I_STAGE_LUT[1458] = -16'd201;
assign W_R_STAGE_LUT[1459] = -16'd158;
assign W_I_STAGE_LUT[1459] = -16'd201;
assign W_R_STAGE_LUT[1460] = -16'd159;
assign W_I_STAGE_LUT[1460] = -16'd201;
assign W_R_STAGE_LUT[1461] = -16'd159;
assign W_I_STAGE_LUT[1461] = -16'd201;
assign W_R_STAGE_LUT[1462] = -16'd159;
assign W_I_STAGE_LUT[1462] = -16'd200;
assign W_R_STAGE_LUT[1463] = -16'd160;
assign W_I_STAGE_LUT[1463] = -16'd200;
assign W_R_STAGE_LUT[1464] = -16'd160;
assign W_I_STAGE_LUT[1464] = -16'd200;
assign W_R_STAGE_LUT[1465] = -16'd160;
assign W_I_STAGE_LUT[1465] = -16'd200;
assign W_R_STAGE_LUT[1466] = -16'd161;
assign W_I_STAGE_LUT[1466] = -16'd199;
assign W_R_STAGE_LUT[1467] = -16'd161;
assign W_I_STAGE_LUT[1467] = -16'd199;
assign W_R_STAGE_LUT[1468] = -16'd161;
assign W_I_STAGE_LUT[1468] = -16'd199;
assign W_R_STAGE_LUT[1469] = -16'd161;
assign W_I_STAGE_LUT[1469] = -16'd199;
assign W_R_STAGE_LUT[1470] = -16'd162;
assign W_I_STAGE_LUT[1470] = -16'd198;
assign W_R_STAGE_LUT[1471] = -16'd162;
assign W_I_STAGE_LUT[1471] = -16'd198;
assign W_R_STAGE_LUT[1472] = -16'd162;
assign W_I_STAGE_LUT[1472] = -16'd198;
assign W_R_STAGE_LUT[1473] = -16'd163;
assign W_I_STAGE_LUT[1473] = -16'd198;
assign W_R_STAGE_LUT[1474] = -16'd163;
assign W_I_STAGE_LUT[1474] = -16'd197;
assign W_R_STAGE_LUT[1475] = -16'd163;
assign W_I_STAGE_LUT[1475] = -16'd197;
assign W_R_STAGE_LUT[1476] = -16'd164;
assign W_I_STAGE_LUT[1476] = -16'd197;
assign W_R_STAGE_LUT[1477] = -16'd164;
assign W_I_STAGE_LUT[1477] = -16'd197;
assign W_R_STAGE_LUT[1478] = -16'd164;
assign W_I_STAGE_LUT[1478] = -16'd196;
assign W_R_STAGE_LUT[1479] = -16'd165;
assign W_I_STAGE_LUT[1479] = -16'd196;
assign W_R_STAGE_LUT[1480] = -16'd165;
assign W_I_STAGE_LUT[1480] = -16'd196;
assign W_R_STAGE_LUT[1481] = -16'd165;
assign W_I_STAGE_LUT[1481] = -16'd196;
assign W_R_STAGE_LUT[1482] = -16'd165;
assign W_I_STAGE_LUT[1482] = -16'd195;
assign W_R_STAGE_LUT[1483] = -16'd166;
assign W_I_STAGE_LUT[1483] = -16'd195;
assign W_R_STAGE_LUT[1484] = -16'd166;
assign W_I_STAGE_LUT[1484] = -16'd195;
assign W_R_STAGE_LUT[1485] = -16'd166;
assign W_I_STAGE_LUT[1485] = -16'd195;
assign W_R_STAGE_LUT[1486] = -16'd167;
assign W_I_STAGE_LUT[1486] = -16'd194;
assign W_R_STAGE_LUT[1487] = -16'd167;
assign W_I_STAGE_LUT[1487] = -16'd194;
assign W_R_STAGE_LUT[1488] = -16'd167;
assign W_I_STAGE_LUT[1488] = -16'd194;
assign W_R_STAGE_LUT[1489] = -16'd168;
assign W_I_STAGE_LUT[1489] = -16'd194;
assign W_R_STAGE_LUT[1490] = -16'd168;
assign W_I_STAGE_LUT[1490] = -16'd193;
assign W_R_STAGE_LUT[1491] = -16'd168;
assign W_I_STAGE_LUT[1491] = -16'd193;
assign W_R_STAGE_LUT[1492] = -16'd168;
assign W_I_STAGE_LUT[1492] = -16'd193;
assign W_R_STAGE_LUT[1493] = -16'd169;
assign W_I_STAGE_LUT[1493] = -16'd193;
assign W_R_STAGE_LUT[1494] = -16'd169;
assign W_I_STAGE_LUT[1494] = -16'd192;
assign W_R_STAGE_LUT[1495] = -16'd169;
assign W_I_STAGE_LUT[1495] = -16'd192;
assign W_R_STAGE_LUT[1496] = -16'd170;
assign W_I_STAGE_LUT[1496] = -16'd192;
assign W_R_STAGE_LUT[1497] = -16'd170;
assign W_I_STAGE_LUT[1497] = -16'd192;
assign W_R_STAGE_LUT[1498] = -16'd170;
assign W_I_STAGE_LUT[1498] = -16'd191;
assign W_R_STAGE_LUT[1499] = -16'd170;
assign W_I_STAGE_LUT[1499] = -16'd191;
assign W_R_STAGE_LUT[1500] = -16'd171;
assign W_I_STAGE_LUT[1500] = -16'd191;
assign W_R_STAGE_LUT[1501] = -16'd171;
assign W_I_STAGE_LUT[1501] = -16'd190;
assign W_R_STAGE_LUT[1502] = -16'd171;
assign W_I_STAGE_LUT[1502] = -16'd190;
assign W_R_STAGE_LUT[1503] = -16'd172;
assign W_I_STAGE_LUT[1503] = -16'd190;
assign W_R_STAGE_LUT[1504] = -16'd172;
assign W_I_STAGE_LUT[1504] = -16'd190;
assign W_R_STAGE_LUT[1505] = -16'd172;
assign W_I_STAGE_LUT[1505] = -16'd189;
assign W_R_STAGE_LUT[1506] = -16'd173;
assign W_I_STAGE_LUT[1506] = -16'd189;
assign W_R_STAGE_LUT[1507] = -16'd173;
assign W_I_STAGE_LUT[1507] = -16'd189;
assign W_R_STAGE_LUT[1508] = -16'd173;
assign W_I_STAGE_LUT[1508] = -16'd189;
assign W_R_STAGE_LUT[1509] = -16'd173;
assign W_I_STAGE_LUT[1509] = -16'd188;
assign W_R_STAGE_LUT[1510] = -16'd174;
assign W_I_STAGE_LUT[1510] = -16'd188;
assign W_R_STAGE_LUT[1511] = -16'd174;
assign W_I_STAGE_LUT[1511] = -16'd188;
assign W_R_STAGE_LUT[1512] = -16'd174;
assign W_I_STAGE_LUT[1512] = -16'd188;
assign W_R_STAGE_LUT[1513] = -16'd175;
assign W_I_STAGE_LUT[1513] = -16'd187;
assign W_R_STAGE_LUT[1514] = -16'd175;
assign W_I_STAGE_LUT[1514] = -16'd187;
assign W_R_STAGE_LUT[1515] = -16'd175;
assign W_I_STAGE_LUT[1515] = -16'd187;
assign W_R_STAGE_LUT[1516] = -16'd175;
assign W_I_STAGE_LUT[1516] = -16'd186;
assign W_R_STAGE_LUT[1517] = -16'd176;
assign W_I_STAGE_LUT[1517] = -16'd186;
assign W_R_STAGE_LUT[1518] = -16'd176;
assign W_I_STAGE_LUT[1518] = -16'd186;
assign W_R_STAGE_LUT[1519] = -16'd176;
assign W_I_STAGE_LUT[1519] = -16'd186;
assign W_R_STAGE_LUT[1520] = -16'd177;
assign W_I_STAGE_LUT[1520] = -16'd185;
assign W_R_STAGE_LUT[1521] = -16'd177;
assign W_I_STAGE_LUT[1521] = -16'd185;
assign W_R_STAGE_LUT[1522] = -16'd177;
assign W_I_STAGE_LUT[1522] = -16'd185;
assign W_R_STAGE_LUT[1523] = -16'd177;
assign W_I_STAGE_LUT[1523] = -16'd185;
assign W_R_STAGE_LUT[1524] = -16'd178;
assign W_I_STAGE_LUT[1524] = -16'd184;
assign W_R_STAGE_LUT[1525] = -16'd178;
assign W_I_STAGE_LUT[1525] = -16'd184;
assign W_R_STAGE_LUT[1526] = -16'd178;
assign W_I_STAGE_LUT[1526] = -16'd184;
assign W_R_STAGE_LUT[1527] = -16'd179;
assign W_I_STAGE_LUT[1527] = -16'd184;
assign W_R_STAGE_LUT[1528] = -16'd179;
assign W_I_STAGE_LUT[1528] = -16'd183;
assign W_R_STAGE_LUT[1529] = -16'd179;
assign W_I_STAGE_LUT[1529] = -16'd183;
assign W_R_STAGE_LUT[1530] = -16'd179;
assign W_I_STAGE_LUT[1530] = -16'd183;
assign W_R_STAGE_LUT[1531] = -16'd180;
assign W_I_STAGE_LUT[1531] = -16'd182;
assign W_R_STAGE_LUT[1532] = -16'd180;
assign W_I_STAGE_LUT[1532] = -16'd182;
assign W_R_STAGE_LUT[1533] = -16'd180;
assign W_I_STAGE_LUT[1533] = -16'd182;
assign W_R_STAGE_LUT[1534] = -16'd180;
assign W_I_STAGE_LUT[1534] = -16'd182;
assign W_R_STAGE_LUT[1535] = -16'd181;
assign W_I_STAGE_LUT[1535] = -16'd181;
assign W_R_STAGE_LUT[1536] = -16'd181;
assign W_I_STAGE_LUT[1536] = -16'd181;
assign W_R_STAGE_LUT[1537] = -16'd181;
assign W_I_STAGE_LUT[1537] = -16'd181;
assign W_R_STAGE_LUT[1538] = -16'd182;
assign W_I_STAGE_LUT[1538] = -16'd180;
assign W_R_STAGE_LUT[1539] = -16'd182;
assign W_I_STAGE_LUT[1539] = -16'd180;
assign W_R_STAGE_LUT[1540] = -16'd182;
assign W_I_STAGE_LUT[1540] = -16'd180;
assign W_R_STAGE_LUT[1541] = -16'd182;
assign W_I_STAGE_LUT[1541] = -16'd180;
assign W_R_STAGE_LUT[1542] = -16'd183;
assign W_I_STAGE_LUT[1542] = -16'd179;
assign W_R_STAGE_LUT[1543] = -16'd183;
assign W_I_STAGE_LUT[1543] = -16'd179;
assign W_R_STAGE_LUT[1544] = -16'd183;
assign W_I_STAGE_LUT[1544] = -16'd179;
assign W_R_STAGE_LUT[1545] = -16'd184;
assign W_I_STAGE_LUT[1545] = -16'd179;
assign W_R_STAGE_LUT[1546] = -16'd184;
assign W_I_STAGE_LUT[1546] = -16'd178;
assign W_R_STAGE_LUT[1547] = -16'd184;
assign W_I_STAGE_LUT[1547] = -16'd178;
assign W_R_STAGE_LUT[1548] = -16'd184;
assign W_I_STAGE_LUT[1548] = -16'd178;
assign W_R_STAGE_LUT[1549] = -16'd185;
assign W_I_STAGE_LUT[1549] = -16'd177;
assign W_R_STAGE_LUT[1550] = -16'd185;
assign W_I_STAGE_LUT[1550] = -16'd177;
assign W_R_STAGE_LUT[1551] = -16'd185;
assign W_I_STAGE_LUT[1551] = -16'd177;
assign W_R_STAGE_LUT[1552] = -16'd185;
assign W_I_STAGE_LUT[1552] = -16'd177;
assign W_R_STAGE_LUT[1553] = -16'd186;
assign W_I_STAGE_LUT[1553] = -16'd176;
assign W_R_STAGE_LUT[1554] = -16'd186;
assign W_I_STAGE_LUT[1554] = -16'd176;
assign W_R_STAGE_LUT[1555] = -16'd186;
assign W_I_STAGE_LUT[1555] = -16'd176;
assign W_R_STAGE_LUT[1556] = -16'd186;
assign W_I_STAGE_LUT[1556] = -16'd175;
assign W_R_STAGE_LUT[1557] = -16'd187;
assign W_I_STAGE_LUT[1557] = -16'd175;
assign W_R_STAGE_LUT[1558] = -16'd187;
assign W_I_STAGE_LUT[1558] = -16'd175;
assign W_R_STAGE_LUT[1559] = -16'd187;
assign W_I_STAGE_LUT[1559] = -16'd175;
assign W_R_STAGE_LUT[1560] = -16'd188;
assign W_I_STAGE_LUT[1560] = -16'd174;
assign W_R_STAGE_LUT[1561] = -16'd188;
assign W_I_STAGE_LUT[1561] = -16'd174;
assign W_R_STAGE_LUT[1562] = -16'd188;
assign W_I_STAGE_LUT[1562] = -16'd174;
assign W_R_STAGE_LUT[1563] = -16'd188;
assign W_I_STAGE_LUT[1563] = -16'd173;
assign W_R_STAGE_LUT[1564] = -16'd189;
assign W_I_STAGE_LUT[1564] = -16'd173;
assign W_R_STAGE_LUT[1565] = -16'd189;
assign W_I_STAGE_LUT[1565] = -16'd173;
assign W_R_STAGE_LUT[1566] = -16'd189;
assign W_I_STAGE_LUT[1566] = -16'd173;
assign W_R_STAGE_LUT[1567] = -16'd189;
assign W_I_STAGE_LUT[1567] = -16'd172;
assign W_R_STAGE_LUT[1568] = -16'd190;
assign W_I_STAGE_LUT[1568] = -16'd172;
assign W_R_STAGE_LUT[1569] = -16'd190;
assign W_I_STAGE_LUT[1569] = -16'd172;
assign W_R_STAGE_LUT[1570] = -16'd190;
assign W_I_STAGE_LUT[1570] = -16'd171;
assign W_R_STAGE_LUT[1571] = -16'd190;
assign W_I_STAGE_LUT[1571] = -16'd171;
assign W_R_STAGE_LUT[1572] = -16'd191;
assign W_I_STAGE_LUT[1572] = -16'd171;
assign W_R_STAGE_LUT[1573] = -16'd191;
assign W_I_STAGE_LUT[1573] = -16'd170;
assign W_R_STAGE_LUT[1574] = -16'd191;
assign W_I_STAGE_LUT[1574] = -16'd170;
assign W_R_STAGE_LUT[1575] = -16'd192;
assign W_I_STAGE_LUT[1575] = -16'd170;
assign W_R_STAGE_LUT[1576] = -16'd192;
assign W_I_STAGE_LUT[1576] = -16'd170;
assign W_R_STAGE_LUT[1577] = -16'd192;
assign W_I_STAGE_LUT[1577] = -16'd169;
assign W_R_STAGE_LUT[1578] = -16'd192;
assign W_I_STAGE_LUT[1578] = -16'd169;
assign W_R_STAGE_LUT[1579] = -16'd193;
assign W_I_STAGE_LUT[1579] = -16'd169;
assign W_R_STAGE_LUT[1580] = -16'd193;
assign W_I_STAGE_LUT[1580] = -16'd168;
assign W_R_STAGE_LUT[1581] = -16'd193;
assign W_I_STAGE_LUT[1581] = -16'd168;
assign W_R_STAGE_LUT[1582] = -16'd193;
assign W_I_STAGE_LUT[1582] = -16'd168;
assign W_R_STAGE_LUT[1583] = -16'd194;
assign W_I_STAGE_LUT[1583] = -16'd168;
assign W_R_STAGE_LUT[1584] = -16'd194;
assign W_I_STAGE_LUT[1584] = -16'd167;
assign W_R_STAGE_LUT[1585] = -16'd194;
assign W_I_STAGE_LUT[1585] = -16'd167;
assign W_R_STAGE_LUT[1586] = -16'd194;
assign W_I_STAGE_LUT[1586] = -16'd167;
assign W_R_STAGE_LUT[1587] = -16'd195;
assign W_I_STAGE_LUT[1587] = -16'd166;
assign W_R_STAGE_LUT[1588] = -16'd195;
assign W_I_STAGE_LUT[1588] = -16'd166;
assign W_R_STAGE_LUT[1589] = -16'd195;
assign W_I_STAGE_LUT[1589] = -16'd166;
assign W_R_STAGE_LUT[1590] = -16'd195;
assign W_I_STAGE_LUT[1590] = -16'd165;
assign W_R_STAGE_LUT[1591] = -16'd196;
assign W_I_STAGE_LUT[1591] = -16'd165;
assign W_R_STAGE_LUT[1592] = -16'd196;
assign W_I_STAGE_LUT[1592] = -16'd165;
assign W_R_STAGE_LUT[1593] = -16'd196;
assign W_I_STAGE_LUT[1593] = -16'd165;
assign W_R_STAGE_LUT[1594] = -16'd196;
assign W_I_STAGE_LUT[1594] = -16'd164;
assign W_R_STAGE_LUT[1595] = -16'd197;
assign W_I_STAGE_LUT[1595] = -16'd164;
assign W_R_STAGE_LUT[1596] = -16'd197;
assign W_I_STAGE_LUT[1596] = -16'd164;
assign W_R_STAGE_LUT[1597] = -16'd197;
assign W_I_STAGE_LUT[1597] = -16'd163;
assign W_R_STAGE_LUT[1598] = -16'd197;
assign W_I_STAGE_LUT[1598] = -16'd163;
assign W_R_STAGE_LUT[1599] = -16'd198;
assign W_I_STAGE_LUT[1599] = -16'd163;
assign W_R_STAGE_LUT[1600] = -16'd198;
assign W_I_STAGE_LUT[1600] = -16'd162;
assign W_R_STAGE_LUT[1601] = -16'd198;
assign W_I_STAGE_LUT[1601] = -16'd162;
assign W_R_STAGE_LUT[1602] = -16'd198;
assign W_I_STAGE_LUT[1602] = -16'd162;
assign W_R_STAGE_LUT[1603] = -16'd199;
assign W_I_STAGE_LUT[1603] = -16'd161;
assign W_R_STAGE_LUT[1604] = -16'd199;
assign W_I_STAGE_LUT[1604] = -16'd161;
assign W_R_STAGE_LUT[1605] = -16'd199;
assign W_I_STAGE_LUT[1605] = -16'd161;
assign W_R_STAGE_LUT[1606] = -16'd199;
assign W_I_STAGE_LUT[1606] = -16'd161;
assign W_R_STAGE_LUT[1607] = -16'd200;
assign W_I_STAGE_LUT[1607] = -16'd160;
assign W_R_STAGE_LUT[1608] = -16'd200;
assign W_I_STAGE_LUT[1608] = -16'd160;
assign W_R_STAGE_LUT[1609] = -16'd200;
assign W_I_STAGE_LUT[1609] = -16'd160;
assign W_R_STAGE_LUT[1610] = -16'd200;
assign W_I_STAGE_LUT[1610] = -16'd159;
assign W_R_STAGE_LUT[1611] = -16'd201;
assign W_I_STAGE_LUT[1611] = -16'd159;
assign W_R_STAGE_LUT[1612] = -16'd201;
assign W_I_STAGE_LUT[1612] = -16'd159;
assign W_R_STAGE_LUT[1613] = -16'd201;
assign W_I_STAGE_LUT[1613] = -16'd158;
assign W_R_STAGE_LUT[1614] = -16'd201;
assign W_I_STAGE_LUT[1614] = -16'd158;
assign W_R_STAGE_LUT[1615] = -16'd202;
assign W_I_STAGE_LUT[1615] = -16'd158;
assign W_R_STAGE_LUT[1616] = -16'd202;
assign W_I_STAGE_LUT[1616] = -16'd157;
assign W_R_STAGE_LUT[1617] = -16'd202;
assign W_I_STAGE_LUT[1617] = -16'd157;
assign W_R_STAGE_LUT[1618] = -16'd202;
assign W_I_STAGE_LUT[1618] = -16'd157;
assign W_R_STAGE_LUT[1619] = -16'd203;
assign W_I_STAGE_LUT[1619] = -16'd157;
assign W_R_STAGE_LUT[1620] = -16'd203;
assign W_I_STAGE_LUT[1620] = -16'd156;
assign W_R_STAGE_LUT[1621] = -16'd203;
assign W_I_STAGE_LUT[1621] = -16'd156;
assign W_R_STAGE_LUT[1622] = -16'd203;
assign W_I_STAGE_LUT[1622] = -16'd156;
assign W_R_STAGE_LUT[1623] = -16'd203;
assign W_I_STAGE_LUT[1623] = -16'd155;
assign W_R_STAGE_LUT[1624] = -16'd204;
assign W_I_STAGE_LUT[1624] = -16'd155;
assign W_R_STAGE_LUT[1625] = -16'd204;
assign W_I_STAGE_LUT[1625] = -16'd155;
assign W_R_STAGE_LUT[1626] = -16'd204;
assign W_I_STAGE_LUT[1626] = -16'd154;
assign W_R_STAGE_LUT[1627] = -16'd204;
assign W_I_STAGE_LUT[1627] = -16'd154;
assign W_R_STAGE_LUT[1628] = -16'd205;
assign W_I_STAGE_LUT[1628] = -16'd154;
assign W_R_STAGE_LUT[1629] = -16'd205;
assign W_I_STAGE_LUT[1629] = -16'd153;
assign W_R_STAGE_LUT[1630] = -16'd205;
assign W_I_STAGE_LUT[1630] = -16'd153;
assign W_R_STAGE_LUT[1631] = -16'd205;
assign W_I_STAGE_LUT[1631] = -16'd153;
assign W_R_STAGE_LUT[1632] = -16'd206;
assign W_I_STAGE_LUT[1632] = -16'd152;
assign W_R_STAGE_LUT[1633] = -16'd206;
assign W_I_STAGE_LUT[1633] = -16'd152;
assign W_R_STAGE_LUT[1634] = -16'd206;
assign W_I_STAGE_LUT[1634] = -16'd152;
assign W_R_STAGE_LUT[1635] = -16'd206;
assign W_I_STAGE_LUT[1635] = -16'd152;
assign W_R_STAGE_LUT[1636] = -16'd207;
assign W_I_STAGE_LUT[1636] = -16'd151;
assign W_R_STAGE_LUT[1637] = -16'd207;
assign W_I_STAGE_LUT[1637] = -16'd151;
assign W_R_STAGE_LUT[1638] = -16'd207;
assign W_I_STAGE_LUT[1638] = -16'd151;
assign W_R_STAGE_LUT[1639] = -16'd207;
assign W_I_STAGE_LUT[1639] = -16'd150;
assign W_R_STAGE_LUT[1640] = -16'd207;
assign W_I_STAGE_LUT[1640] = -16'd150;
assign W_R_STAGE_LUT[1641] = -16'd208;
assign W_I_STAGE_LUT[1641] = -16'd150;
assign W_R_STAGE_LUT[1642] = -16'd208;
assign W_I_STAGE_LUT[1642] = -16'd149;
assign W_R_STAGE_LUT[1643] = -16'd208;
assign W_I_STAGE_LUT[1643] = -16'd149;
assign W_R_STAGE_LUT[1644] = -16'd208;
assign W_I_STAGE_LUT[1644] = -16'd149;
assign W_R_STAGE_LUT[1645] = -16'd209;
assign W_I_STAGE_LUT[1645] = -16'd148;
assign W_R_STAGE_LUT[1646] = -16'd209;
assign W_I_STAGE_LUT[1646] = -16'd148;
assign W_R_STAGE_LUT[1647] = -16'd209;
assign W_I_STAGE_LUT[1647] = -16'd148;
assign W_R_STAGE_LUT[1648] = -16'd209;
assign W_I_STAGE_LUT[1648] = -16'd147;
assign W_R_STAGE_LUT[1649] = -16'd210;
assign W_I_STAGE_LUT[1649] = -16'd147;
assign W_R_STAGE_LUT[1650] = -16'd210;
assign W_I_STAGE_LUT[1650] = -16'd147;
assign W_R_STAGE_LUT[1651] = -16'd210;
assign W_I_STAGE_LUT[1651] = -16'd146;
assign W_R_STAGE_LUT[1652] = -16'd210;
assign W_I_STAGE_LUT[1652] = -16'd146;
assign W_R_STAGE_LUT[1653] = -16'd210;
assign W_I_STAGE_LUT[1653] = -16'd146;
assign W_R_STAGE_LUT[1654] = -16'd211;
assign W_I_STAGE_LUT[1654] = -16'd145;
assign W_R_STAGE_LUT[1655] = -16'd211;
assign W_I_STAGE_LUT[1655] = -16'd145;
assign W_R_STAGE_LUT[1656] = -16'd211;
assign W_I_STAGE_LUT[1656] = -16'd145;
assign W_R_STAGE_LUT[1657] = -16'd211;
assign W_I_STAGE_LUT[1657] = -16'd145;
assign W_R_STAGE_LUT[1658] = -16'd212;
assign W_I_STAGE_LUT[1658] = -16'd144;
assign W_R_STAGE_LUT[1659] = -16'd212;
assign W_I_STAGE_LUT[1659] = -16'd144;
assign W_R_STAGE_LUT[1660] = -16'd212;
assign W_I_STAGE_LUT[1660] = -16'd144;
assign W_R_STAGE_LUT[1661] = -16'd212;
assign W_I_STAGE_LUT[1661] = -16'd143;
assign W_R_STAGE_LUT[1662] = -16'd212;
assign W_I_STAGE_LUT[1662] = -16'd143;
assign W_R_STAGE_LUT[1663] = -16'd213;
assign W_I_STAGE_LUT[1663] = -16'd143;
assign W_R_STAGE_LUT[1664] = -16'd213;
assign W_I_STAGE_LUT[1664] = -16'd142;
assign W_R_STAGE_LUT[1665] = -16'd213;
assign W_I_STAGE_LUT[1665] = -16'd142;
assign W_R_STAGE_LUT[1666] = -16'd213;
assign W_I_STAGE_LUT[1666] = -16'd142;
assign W_R_STAGE_LUT[1667] = -16'd214;
assign W_I_STAGE_LUT[1667] = -16'd141;
assign W_R_STAGE_LUT[1668] = -16'd214;
assign W_I_STAGE_LUT[1668] = -16'd141;
assign W_R_STAGE_LUT[1669] = -16'd214;
assign W_I_STAGE_LUT[1669] = -16'd141;
assign W_R_STAGE_LUT[1670] = -16'd214;
assign W_I_STAGE_LUT[1670] = -16'd140;
assign W_R_STAGE_LUT[1671] = -16'd214;
assign W_I_STAGE_LUT[1671] = -16'd140;
assign W_R_STAGE_LUT[1672] = -16'd215;
assign W_I_STAGE_LUT[1672] = -16'd140;
assign W_R_STAGE_LUT[1673] = -16'd215;
assign W_I_STAGE_LUT[1673] = -16'd139;
assign W_R_STAGE_LUT[1674] = -16'd215;
assign W_I_STAGE_LUT[1674] = -16'd139;
assign W_R_STAGE_LUT[1675] = -16'd215;
assign W_I_STAGE_LUT[1675] = -16'd139;
assign W_R_STAGE_LUT[1676] = -16'd215;
assign W_I_STAGE_LUT[1676] = -16'd138;
assign W_R_STAGE_LUT[1677] = -16'd216;
assign W_I_STAGE_LUT[1677] = -16'd138;
assign W_R_STAGE_LUT[1678] = -16'd216;
assign W_I_STAGE_LUT[1678] = -16'd138;
assign W_R_STAGE_LUT[1679] = -16'd216;
assign W_I_STAGE_LUT[1679] = -16'd137;
assign W_R_STAGE_LUT[1680] = -16'd216;
assign W_I_STAGE_LUT[1680] = -16'd137;
assign W_R_STAGE_LUT[1681] = -16'd216;
assign W_I_STAGE_LUT[1681] = -16'd137;
assign W_R_STAGE_LUT[1682] = -16'd217;
assign W_I_STAGE_LUT[1682] = -16'd136;
assign W_R_STAGE_LUT[1683] = -16'd217;
assign W_I_STAGE_LUT[1683] = -16'd136;
assign W_R_STAGE_LUT[1684] = -16'd217;
assign W_I_STAGE_LUT[1684] = -16'd136;
assign W_R_STAGE_LUT[1685] = -16'd217;
assign W_I_STAGE_LUT[1685] = -16'd135;
assign W_R_STAGE_LUT[1686] = -16'd218;
assign W_I_STAGE_LUT[1686] = -16'd135;
assign W_R_STAGE_LUT[1687] = -16'd218;
assign W_I_STAGE_LUT[1687] = -16'd135;
assign W_R_STAGE_LUT[1688] = -16'd218;
assign W_I_STAGE_LUT[1688] = -16'd134;
assign W_R_STAGE_LUT[1689] = -16'd218;
assign W_I_STAGE_LUT[1689] = -16'd134;
assign W_R_STAGE_LUT[1690] = -16'd218;
assign W_I_STAGE_LUT[1690] = -16'd134;
assign W_R_STAGE_LUT[1691] = -16'd219;
assign W_I_STAGE_LUT[1691] = -16'd133;
assign W_R_STAGE_LUT[1692] = -16'd219;
assign W_I_STAGE_LUT[1692] = -16'd133;
assign W_R_STAGE_LUT[1693] = -16'd219;
assign W_I_STAGE_LUT[1693] = -16'd133;
assign W_R_STAGE_LUT[1694] = -16'd219;
assign W_I_STAGE_LUT[1694] = -16'd132;
assign W_R_STAGE_LUT[1695] = -16'd219;
assign W_I_STAGE_LUT[1695] = -16'd132;
assign W_R_STAGE_LUT[1696] = -16'd220;
assign W_I_STAGE_LUT[1696] = -16'd132;
assign W_R_STAGE_LUT[1697] = -16'd220;
assign W_I_STAGE_LUT[1697] = -16'd131;
assign W_R_STAGE_LUT[1698] = -16'd220;
assign W_I_STAGE_LUT[1698] = -16'd131;
assign W_R_STAGE_LUT[1699] = -16'd220;
assign W_I_STAGE_LUT[1699] = -16'd131;
assign W_R_STAGE_LUT[1700] = -16'd220;
assign W_I_STAGE_LUT[1700] = -16'd130;
assign W_R_STAGE_LUT[1701] = -16'd221;
assign W_I_STAGE_LUT[1701] = -16'd130;
assign W_R_STAGE_LUT[1702] = -16'd221;
assign W_I_STAGE_LUT[1702] = -16'd130;
assign W_R_STAGE_LUT[1703] = -16'd221;
assign W_I_STAGE_LUT[1703] = -16'd129;
assign W_R_STAGE_LUT[1704] = -16'd221;
assign W_I_STAGE_LUT[1704] = -16'd129;
assign W_R_STAGE_LUT[1705] = -16'd221;
assign W_I_STAGE_LUT[1705] = -16'd129;
assign W_R_STAGE_LUT[1706] = -16'd222;
assign W_I_STAGE_LUT[1706] = -16'd128;
assign W_R_STAGE_LUT[1707] = -16'd222;
assign W_I_STAGE_LUT[1707] = -16'd128;
assign W_R_STAGE_LUT[1708] = -16'd222;
assign W_I_STAGE_LUT[1708] = -16'd128;
assign W_R_STAGE_LUT[1709] = -16'd222;
assign W_I_STAGE_LUT[1709] = -16'd127;
assign W_R_STAGE_LUT[1710] = -16'd222;
assign W_I_STAGE_LUT[1710] = -16'd127;
assign W_R_STAGE_LUT[1711] = -16'd223;
assign W_I_STAGE_LUT[1711] = -16'd127;
assign W_R_STAGE_LUT[1712] = -16'd223;
assign W_I_STAGE_LUT[1712] = -16'd126;
assign W_R_STAGE_LUT[1713] = -16'd223;
assign W_I_STAGE_LUT[1713] = -16'd126;
assign W_R_STAGE_LUT[1714] = -16'd223;
assign W_I_STAGE_LUT[1714] = -16'd125;
assign W_R_STAGE_LUT[1715] = -16'd223;
assign W_I_STAGE_LUT[1715] = -16'd125;
assign W_R_STAGE_LUT[1716] = -16'd224;
assign W_I_STAGE_LUT[1716] = -16'd125;
assign W_R_STAGE_LUT[1717] = -16'd224;
assign W_I_STAGE_LUT[1717] = -16'd124;
assign W_R_STAGE_LUT[1718] = -16'd224;
assign W_I_STAGE_LUT[1718] = -16'd124;
assign W_R_STAGE_LUT[1719] = -16'd224;
assign W_I_STAGE_LUT[1719] = -16'd124;
assign W_R_STAGE_LUT[1720] = -16'd224;
assign W_I_STAGE_LUT[1720] = -16'd123;
assign W_R_STAGE_LUT[1721] = -16'd224;
assign W_I_STAGE_LUT[1721] = -16'd123;
assign W_R_STAGE_LUT[1722] = -16'd225;
assign W_I_STAGE_LUT[1722] = -16'd123;
assign W_R_STAGE_LUT[1723] = -16'd225;
assign W_I_STAGE_LUT[1723] = -16'd122;
assign W_R_STAGE_LUT[1724] = -16'd225;
assign W_I_STAGE_LUT[1724] = -16'd122;
assign W_R_STAGE_LUT[1725] = -16'd225;
assign W_I_STAGE_LUT[1725] = -16'd122;
assign W_R_STAGE_LUT[1726] = -16'd225;
assign W_I_STAGE_LUT[1726] = -16'd121;
assign W_R_STAGE_LUT[1727] = -16'd226;
assign W_I_STAGE_LUT[1727] = -16'd121;
assign W_R_STAGE_LUT[1728] = -16'd226;
assign W_I_STAGE_LUT[1728] = -16'd121;
assign W_R_STAGE_LUT[1729] = -16'd226;
assign W_I_STAGE_LUT[1729] = -16'd120;
assign W_R_STAGE_LUT[1730] = -16'd226;
assign W_I_STAGE_LUT[1730] = -16'd120;
assign W_R_STAGE_LUT[1731] = -16'd226;
assign W_I_STAGE_LUT[1731] = -16'd120;
assign W_R_STAGE_LUT[1732] = -16'd227;
assign W_I_STAGE_LUT[1732] = -16'd119;
assign W_R_STAGE_LUT[1733] = -16'd227;
assign W_I_STAGE_LUT[1733] = -16'd119;
assign W_R_STAGE_LUT[1734] = -16'd227;
assign W_I_STAGE_LUT[1734] = -16'd119;
assign W_R_STAGE_LUT[1735] = -16'd227;
assign W_I_STAGE_LUT[1735] = -16'd118;
assign W_R_STAGE_LUT[1736] = -16'd227;
assign W_I_STAGE_LUT[1736] = -16'd118;
assign W_R_STAGE_LUT[1737] = -16'd227;
assign W_I_STAGE_LUT[1737] = -16'd118;
assign W_R_STAGE_LUT[1738] = -16'd228;
assign W_I_STAGE_LUT[1738] = -16'd117;
assign W_R_STAGE_LUT[1739] = -16'd228;
assign W_I_STAGE_LUT[1739] = -16'd117;
assign W_R_STAGE_LUT[1740] = -16'd228;
assign W_I_STAGE_LUT[1740] = -16'd117;
assign W_R_STAGE_LUT[1741] = -16'd228;
assign W_I_STAGE_LUT[1741] = -16'd116;
assign W_R_STAGE_LUT[1742] = -16'd228;
assign W_I_STAGE_LUT[1742] = -16'd116;
assign W_R_STAGE_LUT[1743] = -16'd228;
assign W_I_STAGE_LUT[1743] = -16'd115;
assign W_R_STAGE_LUT[1744] = -16'd229;
assign W_I_STAGE_LUT[1744] = -16'd115;
assign W_R_STAGE_LUT[1745] = -16'd229;
assign W_I_STAGE_LUT[1745] = -16'd115;
assign W_R_STAGE_LUT[1746] = -16'd229;
assign W_I_STAGE_LUT[1746] = -16'd114;
assign W_R_STAGE_LUT[1747] = -16'd229;
assign W_I_STAGE_LUT[1747] = -16'd114;
assign W_R_STAGE_LUT[1748] = -16'd229;
assign W_I_STAGE_LUT[1748] = -16'd114;
assign W_R_STAGE_LUT[1749] = -16'd230;
assign W_I_STAGE_LUT[1749] = -16'd113;
assign W_R_STAGE_LUT[1750] = -16'd230;
assign W_I_STAGE_LUT[1750] = -16'd113;
assign W_R_STAGE_LUT[1751] = -16'd230;
assign W_I_STAGE_LUT[1751] = -16'd113;
assign W_R_STAGE_LUT[1752] = -16'd230;
assign W_I_STAGE_LUT[1752] = -16'd112;
assign W_R_STAGE_LUT[1753] = -16'd230;
assign W_I_STAGE_LUT[1753] = -16'd112;
assign W_R_STAGE_LUT[1754] = -16'd230;
assign W_I_STAGE_LUT[1754] = -16'd112;
assign W_R_STAGE_LUT[1755] = -16'd231;
assign W_I_STAGE_LUT[1755] = -16'd111;
assign W_R_STAGE_LUT[1756] = -16'd231;
assign W_I_STAGE_LUT[1756] = -16'd111;
assign W_R_STAGE_LUT[1757] = -16'd231;
assign W_I_STAGE_LUT[1757] = -16'd111;
assign W_R_STAGE_LUT[1758] = -16'd231;
assign W_I_STAGE_LUT[1758] = -16'd110;
assign W_R_STAGE_LUT[1759] = -16'd231;
assign W_I_STAGE_LUT[1759] = -16'd110;
assign W_R_STAGE_LUT[1760] = -16'd231;
assign W_I_STAGE_LUT[1760] = -16'd109;
assign W_R_STAGE_LUT[1761] = -16'd232;
assign W_I_STAGE_LUT[1761] = -16'd109;
assign W_R_STAGE_LUT[1762] = -16'd232;
assign W_I_STAGE_LUT[1762] = -16'd109;
assign W_R_STAGE_LUT[1763] = -16'd232;
assign W_I_STAGE_LUT[1763] = -16'd108;
assign W_R_STAGE_LUT[1764] = -16'd232;
assign W_I_STAGE_LUT[1764] = -16'd108;
assign W_R_STAGE_LUT[1765] = -16'd232;
assign W_I_STAGE_LUT[1765] = -16'd108;
assign W_R_STAGE_LUT[1766] = -16'd232;
assign W_I_STAGE_LUT[1766] = -16'd107;
assign W_R_STAGE_LUT[1767] = -16'd233;
assign W_I_STAGE_LUT[1767] = -16'd107;
assign W_R_STAGE_LUT[1768] = -16'd233;
assign W_I_STAGE_LUT[1768] = -16'd107;
assign W_R_STAGE_LUT[1769] = -16'd233;
assign W_I_STAGE_LUT[1769] = -16'd106;
assign W_R_STAGE_LUT[1770] = -16'd233;
assign W_I_STAGE_LUT[1770] = -16'd106;
assign W_R_STAGE_LUT[1771] = -16'd233;
assign W_I_STAGE_LUT[1771] = -16'd106;
assign W_R_STAGE_LUT[1772] = -16'd233;
assign W_I_STAGE_LUT[1772] = -16'd105;
assign W_R_STAGE_LUT[1773] = -16'd234;
assign W_I_STAGE_LUT[1773] = -16'd105;
assign W_R_STAGE_LUT[1774] = -16'd234;
assign W_I_STAGE_LUT[1774] = -16'd104;
assign W_R_STAGE_LUT[1775] = -16'd234;
assign W_I_STAGE_LUT[1775] = -16'd104;
assign W_R_STAGE_LUT[1776] = -16'd234;
assign W_I_STAGE_LUT[1776] = -16'd104;
assign W_R_STAGE_LUT[1777] = -16'd234;
assign W_I_STAGE_LUT[1777] = -16'd103;
assign W_R_STAGE_LUT[1778] = -16'd234;
assign W_I_STAGE_LUT[1778] = -16'd103;
assign W_R_STAGE_LUT[1779] = -16'd235;
assign W_I_STAGE_LUT[1779] = -16'd103;
assign W_R_STAGE_LUT[1780] = -16'd235;
assign W_I_STAGE_LUT[1780] = -16'd102;
assign W_R_STAGE_LUT[1781] = -16'd235;
assign W_I_STAGE_LUT[1781] = -16'd102;
assign W_R_STAGE_LUT[1782] = -16'd235;
assign W_I_STAGE_LUT[1782] = -16'd102;
assign W_R_STAGE_LUT[1783] = -16'd235;
assign W_I_STAGE_LUT[1783] = -16'd101;
assign W_R_STAGE_LUT[1784] = -16'd235;
assign W_I_STAGE_LUT[1784] = -16'd101;
assign W_R_STAGE_LUT[1785] = -16'd235;
assign W_I_STAGE_LUT[1785] = -16'd101;
assign W_R_STAGE_LUT[1786] = -16'd236;
assign W_I_STAGE_LUT[1786] = -16'd100;
assign W_R_STAGE_LUT[1787] = -16'd236;
assign W_I_STAGE_LUT[1787] = -16'd100;
assign W_R_STAGE_LUT[1788] = -16'd236;
assign W_I_STAGE_LUT[1788] = -16'd99;
assign W_R_STAGE_LUT[1789] = -16'd236;
assign W_I_STAGE_LUT[1789] = -16'd99;
assign W_R_STAGE_LUT[1790] = -16'd236;
assign W_I_STAGE_LUT[1790] = -16'd99;
assign W_R_STAGE_LUT[1791] = -16'd236;
assign W_I_STAGE_LUT[1791] = -16'd98;
assign W_R_STAGE_LUT[1792] = -16'd237;
assign W_I_STAGE_LUT[1792] = -16'd98;
assign W_R_STAGE_LUT[1793] = -16'd237;
assign W_I_STAGE_LUT[1793] = -16'd98;
assign W_R_STAGE_LUT[1794] = -16'd237;
assign W_I_STAGE_LUT[1794] = -16'd97;
assign W_R_STAGE_LUT[1795] = -16'd237;
assign W_I_STAGE_LUT[1795] = -16'd97;
assign W_R_STAGE_LUT[1796] = -16'd237;
assign W_I_STAGE_LUT[1796] = -16'd97;
assign W_R_STAGE_LUT[1797] = -16'd237;
assign W_I_STAGE_LUT[1797] = -16'd96;
assign W_R_STAGE_LUT[1798] = -16'd237;
assign W_I_STAGE_LUT[1798] = -16'd96;
assign W_R_STAGE_LUT[1799] = -16'd238;
assign W_I_STAGE_LUT[1799] = -16'd95;
assign W_R_STAGE_LUT[1800] = -16'd238;
assign W_I_STAGE_LUT[1800] = -16'd95;
assign W_R_STAGE_LUT[1801] = -16'd238;
assign W_I_STAGE_LUT[1801] = -16'd95;
assign W_R_STAGE_LUT[1802] = -16'd238;
assign W_I_STAGE_LUT[1802] = -16'd94;
assign W_R_STAGE_LUT[1803] = -16'd238;
assign W_I_STAGE_LUT[1803] = -16'd94;
assign W_R_STAGE_LUT[1804] = -16'd238;
assign W_I_STAGE_LUT[1804] = -16'd94;
assign W_R_STAGE_LUT[1805] = -16'd238;
assign W_I_STAGE_LUT[1805] = -16'd93;
assign W_R_STAGE_LUT[1806] = -16'd239;
assign W_I_STAGE_LUT[1806] = -16'd93;
assign W_R_STAGE_LUT[1807] = -16'd239;
assign W_I_STAGE_LUT[1807] = -16'd92;
assign W_R_STAGE_LUT[1808] = -16'd239;
assign W_I_STAGE_LUT[1808] = -16'd92;
assign W_R_STAGE_LUT[1809] = -16'd239;
assign W_I_STAGE_LUT[1809] = -16'd92;
assign W_R_STAGE_LUT[1810] = -16'd239;
assign W_I_STAGE_LUT[1810] = -16'd91;
assign W_R_STAGE_LUT[1811] = -16'd239;
assign W_I_STAGE_LUT[1811] = -16'd91;
assign W_R_STAGE_LUT[1812] = -16'd239;
assign W_I_STAGE_LUT[1812] = -16'd91;
assign W_R_STAGE_LUT[1813] = -16'd240;
assign W_I_STAGE_LUT[1813] = -16'd90;
assign W_R_STAGE_LUT[1814] = -16'd240;
assign W_I_STAGE_LUT[1814] = -16'd90;
assign W_R_STAGE_LUT[1815] = -16'd240;
assign W_I_STAGE_LUT[1815] = -16'd90;
assign W_R_STAGE_LUT[1816] = -16'd240;
assign W_I_STAGE_LUT[1816] = -16'd89;
assign W_R_STAGE_LUT[1817] = -16'd240;
assign W_I_STAGE_LUT[1817] = -16'd89;
assign W_R_STAGE_LUT[1818] = -16'd240;
assign W_I_STAGE_LUT[1818] = -16'd88;
assign W_R_STAGE_LUT[1819] = -16'd240;
assign W_I_STAGE_LUT[1819] = -16'd88;
assign W_R_STAGE_LUT[1820] = -16'd241;
assign W_I_STAGE_LUT[1820] = -16'd88;
assign W_R_STAGE_LUT[1821] = -16'd241;
assign W_I_STAGE_LUT[1821] = -16'd87;
assign W_R_STAGE_LUT[1822] = -16'd241;
assign W_I_STAGE_LUT[1822] = -16'd87;
assign W_R_STAGE_LUT[1823] = -16'd241;
assign W_I_STAGE_LUT[1823] = -16'd87;
assign W_R_STAGE_LUT[1824] = -16'd241;
assign W_I_STAGE_LUT[1824] = -16'd86;
assign W_R_STAGE_LUT[1825] = -16'd241;
assign W_I_STAGE_LUT[1825] = -16'd86;
assign W_R_STAGE_LUT[1826] = -16'd241;
assign W_I_STAGE_LUT[1826] = -16'd86;
assign W_R_STAGE_LUT[1827] = -16'd241;
assign W_I_STAGE_LUT[1827] = -16'd85;
assign W_R_STAGE_LUT[1828] = -16'd242;
assign W_I_STAGE_LUT[1828] = -16'd85;
assign W_R_STAGE_LUT[1829] = -16'd242;
assign W_I_STAGE_LUT[1829] = -16'd84;
assign W_R_STAGE_LUT[1830] = -16'd242;
assign W_I_STAGE_LUT[1830] = -16'd84;
assign W_R_STAGE_LUT[1831] = -16'd242;
assign W_I_STAGE_LUT[1831] = -16'd84;
assign W_R_STAGE_LUT[1832] = -16'd242;
assign W_I_STAGE_LUT[1832] = -16'd83;
assign W_R_STAGE_LUT[1833] = -16'd242;
assign W_I_STAGE_LUT[1833] = -16'd83;
assign W_R_STAGE_LUT[1834] = -16'd242;
assign W_I_STAGE_LUT[1834] = -16'd83;
assign W_R_STAGE_LUT[1835] = -16'd242;
assign W_I_STAGE_LUT[1835] = -16'd82;
assign W_R_STAGE_LUT[1836] = -16'd243;
assign W_I_STAGE_LUT[1836] = -16'd82;
assign W_R_STAGE_LUT[1837] = -16'd243;
assign W_I_STAGE_LUT[1837] = -16'd81;
assign W_R_STAGE_LUT[1838] = -16'd243;
assign W_I_STAGE_LUT[1838] = -16'd81;
assign W_R_STAGE_LUT[1839] = -16'd243;
assign W_I_STAGE_LUT[1839] = -16'd81;
assign W_R_STAGE_LUT[1840] = -16'd243;
assign W_I_STAGE_LUT[1840] = -16'd80;
assign W_R_STAGE_LUT[1841] = -16'd243;
assign W_I_STAGE_LUT[1841] = -16'd80;
assign W_R_STAGE_LUT[1842] = -16'd243;
assign W_I_STAGE_LUT[1842] = -16'd80;
assign W_R_STAGE_LUT[1843] = -16'd243;
assign W_I_STAGE_LUT[1843] = -16'd79;
assign W_R_STAGE_LUT[1844] = -16'd244;
assign W_I_STAGE_LUT[1844] = -16'd79;
assign W_R_STAGE_LUT[1845] = -16'd244;
assign W_I_STAGE_LUT[1845] = -16'd78;
assign W_R_STAGE_LUT[1846] = -16'd244;
assign W_I_STAGE_LUT[1846] = -16'd78;
assign W_R_STAGE_LUT[1847] = -16'd244;
assign W_I_STAGE_LUT[1847] = -16'd78;
assign W_R_STAGE_LUT[1848] = -16'd244;
assign W_I_STAGE_LUT[1848] = -16'd77;
assign W_R_STAGE_LUT[1849] = -16'd244;
assign W_I_STAGE_LUT[1849] = -16'd77;
assign W_R_STAGE_LUT[1850] = -16'd244;
assign W_I_STAGE_LUT[1850] = -16'd77;
assign W_R_STAGE_LUT[1851] = -16'd244;
assign W_I_STAGE_LUT[1851] = -16'd76;
assign W_R_STAGE_LUT[1852] = -16'd245;
assign W_I_STAGE_LUT[1852] = -16'd76;
assign W_R_STAGE_LUT[1853] = -16'd245;
assign W_I_STAGE_LUT[1853] = -16'd75;
assign W_R_STAGE_LUT[1854] = -16'd245;
assign W_I_STAGE_LUT[1854] = -16'd75;
assign W_R_STAGE_LUT[1855] = -16'd245;
assign W_I_STAGE_LUT[1855] = -16'd75;
assign W_R_STAGE_LUT[1856] = -16'd245;
assign W_I_STAGE_LUT[1856] = -16'd74;
assign W_R_STAGE_LUT[1857] = -16'd245;
assign W_I_STAGE_LUT[1857] = -16'd74;
assign W_R_STAGE_LUT[1858] = -16'd245;
assign W_I_STAGE_LUT[1858] = -16'd74;
assign W_R_STAGE_LUT[1859] = -16'd245;
assign W_I_STAGE_LUT[1859] = -16'd73;
assign W_R_STAGE_LUT[1860] = -16'd245;
assign W_I_STAGE_LUT[1860] = -16'd73;
assign W_R_STAGE_LUT[1861] = -16'd246;
assign W_I_STAGE_LUT[1861] = -16'd72;
assign W_R_STAGE_LUT[1862] = -16'd246;
assign W_I_STAGE_LUT[1862] = -16'd72;
assign W_R_STAGE_LUT[1863] = -16'd246;
assign W_I_STAGE_LUT[1863] = -16'd72;
assign W_R_STAGE_LUT[1864] = -16'd246;
assign W_I_STAGE_LUT[1864] = -16'd71;
assign W_R_STAGE_LUT[1865] = -16'd246;
assign W_I_STAGE_LUT[1865] = -16'd71;
assign W_R_STAGE_LUT[1866] = -16'd246;
assign W_I_STAGE_LUT[1866] = -16'd71;
assign W_R_STAGE_LUT[1867] = -16'd246;
assign W_I_STAGE_LUT[1867] = -16'd70;
assign W_R_STAGE_LUT[1868] = -16'd246;
assign W_I_STAGE_LUT[1868] = -16'd70;
assign W_R_STAGE_LUT[1869] = -16'd246;
assign W_I_STAGE_LUT[1869] = -16'd69;
assign W_R_STAGE_LUT[1870] = -16'd247;
assign W_I_STAGE_LUT[1870] = -16'd69;
assign W_R_STAGE_LUT[1871] = -16'd247;
assign W_I_STAGE_LUT[1871] = -16'd69;
assign W_R_STAGE_LUT[1872] = -16'd247;
assign W_I_STAGE_LUT[1872] = -16'd68;
assign W_R_STAGE_LUT[1873] = -16'd247;
assign W_I_STAGE_LUT[1873] = -16'd68;
assign W_R_STAGE_LUT[1874] = -16'd247;
assign W_I_STAGE_LUT[1874] = -16'd68;
assign W_R_STAGE_LUT[1875] = -16'd247;
assign W_I_STAGE_LUT[1875] = -16'd67;
assign W_R_STAGE_LUT[1876] = -16'd247;
assign W_I_STAGE_LUT[1876] = -16'd67;
assign W_R_STAGE_LUT[1877] = -16'd247;
assign W_I_STAGE_LUT[1877] = -16'd66;
assign W_R_STAGE_LUT[1878] = -16'd247;
assign W_I_STAGE_LUT[1878] = -16'd66;
assign W_R_STAGE_LUT[1879] = -16'd247;
assign W_I_STAGE_LUT[1879] = -16'd66;
assign W_R_STAGE_LUT[1880] = -16'd248;
assign W_I_STAGE_LUT[1880] = -16'd65;
assign W_R_STAGE_LUT[1881] = -16'd248;
assign W_I_STAGE_LUT[1881] = -16'd65;
assign W_R_STAGE_LUT[1882] = -16'd248;
assign W_I_STAGE_LUT[1882] = -16'd64;
assign W_R_STAGE_LUT[1883] = -16'd248;
assign W_I_STAGE_LUT[1883] = -16'd64;
assign W_R_STAGE_LUT[1884] = -16'd248;
assign W_I_STAGE_LUT[1884] = -16'd64;
assign W_R_STAGE_LUT[1885] = -16'd248;
assign W_I_STAGE_LUT[1885] = -16'd63;
assign W_R_STAGE_LUT[1886] = -16'd248;
assign W_I_STAGE_LUT[1886] = -16'd63;
assign W_R_STAGE_LUT[1887] = -16'd248;
assign W_I_STAGE_LUT[1887] = -16'd63;
assign W_R_STAGE_LUT[1888] = -16'd248;
assign W_I_STAGE_LUT[1888] = -16'd62;
assign W_R_STAGE_LUT[1889] = -16'd248;
assign W_I_STAGE_LUT[1889] = -16'd62;
assign W_R_STAGE_LUT[1890] = -16'd249;
assign W_I_STAGE_LUT[1890] = -16'd61;
assign W_R_STAGE_LUT[1891] = -16'd249;
assign W_I_STAGE_LUT[1891] = -16'd61;
assign W_R_STAGE_LUT[1892] = -16'd249;
assign W_I_STAGE_LUT[1892] = -16'd61;
assign W_R_STAGE_LUT[1893] = -16'd249;
assign W_I_STAGE_LUT[1893] = -16'd60;
assign W_R_STAGE_LUT[1894] = -16'd249;
assign W_I_STAGE_LUT[1894] = -16'd60;
assign W_R_STAGE_LUT[1895] = -16'd249;
assign W_I_STAGE_LUT[1895] = -16'd60;
assign W_R_STAGE_LUT[1896] = -16'd249;
assign W_I_STAGE_LUT[1896] = -16'd59;
assign W_R_STAGE_LUT[1897] = -16'd249;
assign W_I_STAGE_LUT[1897] = -16'd59;
assign W_R_STAGE_LUT[1898] = -16'd249;
assign W_I_STAGE_LUT[1898] = -16'd58;
assign W_R_STAGE_LUT[1899] = -16'd249;
assign W_I_STAGE_LUT[1899] = -16'd58;
assign W_R_STAGE_LUT[1900] = -16'd249;
assign W_I_STAGE_LUT[1900] = -16'd58;
assign W_R_STAGE_LUT[1901] = -16'd250;
assign W_I_STAGE_LUT[1901] = -16'd57;
assign W_R_STAGE_LUT[1902] = -16'd250;
assign W_I_STAGE_LUT[1902] = -16'd57;
assign W_R_STAGE_LUT[1903] = -16'd250;
assign W_I_STAGE_LUT[1903] = -16'd56;
assign W_R_STAGE_LUT[1904] = -16'd250;
assign W_I_STAGE_LUT[1904] = -16'd56;
assign W_R_STAGE_LUT[1905] = -16'd250;
assign W_I_STAGE_LUT[1905] = -16'd56;
assign W_R_STAGE_LUT[1906] = -16'd250;
assign W_I_STAGE_LUT[1906] = -16'd55;
assign W_R_STAGE_LUT[1907] = -16'd250;
assign W_I_STAGE_LUT[1907] = -16'd55;
assign W_R_STAGE_LUT[1908] = -16'd250;
assign W_I_STAGE_LUT[1908] = -16'd55;
assign W_R_STAGE_LUT[1909] = -16'd250;
assign W_I_STAGE_LUT[1909] = -16'd54;
assign W_R_STAGE_LUT[1910] = -16'd250;
assign W_I_STAGE_LUT[1910] = -16'd54;
assign W_R_STAGE_LUT[1911] = -16'd250;
assign W_I_STAGE_LUT[1911] = -16'd53;
assign W_R_STAGE_LUT[1912] = -16'd250;
assign W_I_STAGE_LUT[1912] = -16'd53;
assign W_R_STAGE_LUT[1913] = -16'd251;
assign W_I_STAGE_LUT[1913] = -16'd53;
assign W_R_STAGE_LUT[1914] = -16'd251;
assign W_I_STAGE_LUT[1914] = -16'd52;
assign W_R_STAGE_LUT[1915] = -16'd251;
assign W_I_STAGE_LUT[1915] = -16'd52;
assign W_R_STAGE_LUT[1916] = -16'd251;
assign W_I_STAGE_LUT[1916] = -16'd51;
assign W_R_STAGE_LUT[1917] = -16'd251;
assign W_I_STAGE_LUT[1917] = -16'd51;
assign W_R_STAGE_LUT[1918] = -16'd251;
assign W_I_STAGE_LUT[1918] = -16'd51;
assign W_R_STAGE_LUT[1919] = -16'd251;
assign W_I_STAGE_LUT[1919] = -16'd50;
assign W_R_STAGE_LUT[1920] = -16'd251;
assign W_I_STAGE_LUT[1920] = -16'd50;
assign W_R_STAGE_LUT[1921] = -16'd251;
assign W_I_STAGE_LUT[1921] = -16'd50;
assign W_R_STAGE_LUT[1922] = -16'd251;
assign W_I_STAGE_LUT[1922] = -16'd49;
assign W_R_STAGE_LUT[1923] = -16'd251;
assign W_I_STAGE_LUT[1923] = -16'd49;
assign W_R_STAGE_LUT[1924] = -16'd251;
assign W_I_STAGE_LUT[1924] = -16'd48;
assign W_R_STAGE_LUT[1925] = -16'd251;
assign W_I_STAGE_LUT[1925] = -16'd48;
assign W_R_STAGE_LUT[1926] = -16'd252;
assign W_I_STAGE_LUT[1926] = -16'd48;
assign W_R_STAGE_LUT[1927] = -16'd252;
assign W_I_STAGE_LUT[1927] = -16'd47;
assign W_R_STAGE_LUT[1928] = -16'd252;
assign W_I_STAGE_LUT[1928] = -16'd47;
assign W_R_STAGE_LUT[1929] = -16'd252;
assign W_I_STAGE_LUT[1929] = -16'd46;
assign W_R_STAGE_LUT[1930] = -16'd252;
assign W_I_STAGE_LUT[1930] = -16'd46;
assign W_R_STAGE_LUT[1931] = -16'd252;
assign W_I_STAGE_LUT[1931] = -16'd46;
assign W_R_STAGE_LUT[1932] = -16'd252;
assign W_I_STAGE_LUT[1932] = -16'd45;
assign W_R_STAGE_LUT[1933] = -16'd252;
assign W_I_STAGE_LUT[1933] = -16'd45;
assign W_R_STAGE_LUT[1934] = -16'd252;
assign W_I_STAGE_LUT[1934] = -16'd45;
assign W_R_STAGE_LUT[1935] = -16'd252;
assign W_I_STAGE_LUT[1935] = -16'd44;
assign W_R_STAGE_LUT[1936] = -16'd252;
assign W_I_STAGE_LUT[1936] = -16'd44;
assign W_R_STAGE_LUT[1937] = -16'd252;
assign W_I_STAGE_LUT[1937] = -16'd43;
assign W_R_STAGE_LUT[1938] = -16'd252;
assign W_I_STAGE_LUT[1938] = -16'd43;
assign W_R_STAGE_LUT[1939] = -16'd252;
assign W_I_STAGE_LUT[1939] = -16'd43;
assign W_R_STAGE_LUT[1940] = -16'd252;
assign W_I_STAGE_LUT[1940] = -16'd42;
assign W_R_STAGE_LUT[1941] = -16'd253;
assign W_I_STAGE_LUT[1941] = -16'd42;
assign W_R_STAGE_LUT[1942] = -16'd253;
assign W_I_STAGE_LUT[1942] = -16'd41;
assign W_R_STAGE_LUT[1943] = -16'd253;
assign W_I_STAGE_LUT[1943] = -16'd41;
assign W_R_STAGE_LUT[1944] = -16'd253;
assign W_I_STAGE_LUT[1944] = -16'd41;
assign W_R_STAGE_LUT[1945] = -16'd253;
assign W_I_STAGE_LUT[1945] = -16'd40;
assign W_R_STAGE_LUT[1946] = -16'd253;
assign W_I_STAGE_LUT[1946] = -16'd40;
assign W_R_STAGE_LUT[1947] = -16'd253;
assign W_I_STAGE_LUT[1947] = -16'd40;
assign W_R_STAGE_LUT[1948] = -16'd253;
assign W_I_STAGE_LUT[1948] = -16'd39;
assign W_R_STAGE_LUT[1949] = -16'd253;
assign W_I_STAGE_LUT[1949] = -16'd39;
assign W_R_STAGE_LUT[1950] = -16'd253;
assign W_I_STAGE_LUT[1950] = -16'd38;
assign W_R_STAGE_LUT[1951] = -16'd253;
assign W_I_STAGE_LUT[1951] = -16'd38;
assign W_R_STAGE_LUT[1952] = -16'd253;
assign W_I_STAGE_LUT[1952] = -16'd38;
assign W_R_STAGE_LUT[1953] = -16'd253;
assign W_I_STAGE_LUT[1953] = -16'd37;
assign W_R_STAGE_LUT[1954] = -16'd253;
assign W_I_STAGE_LUT[1954] = -16'd37;
assign W_R_STAGE_LUT[1955] = -16'd253;
assign W_I_STAGE_LUT[1955] = -16'd36;
assign W_R_STAGE_LUT[1956] = -16'd253;
assign W_I_STAGE_LUT[1956] = -16'd36;
assign W_R_STAGE_LUT[1957] = -16'd254;
assign W_I_STAGE_LUT[1957] = -16'd36;
assign W_R_STAGE_LUT[1958] = -16'd254;
assign W_I_STAGE_LUT[1958] = -16'd35;
assign W_R_STAGE_LUT[1959] = -16'd254;
assign W_I_STAGE_LUT[1959] = -16'd35;
assign W_R_STAGE_LUT[1960] = -16'd254;
assign W_I_STAGE_LUT[1960] = -16'd34;
assign W_R_STAGE_LUT[1961] = -16'd254;
assign W_I_STAGE_LUT[1961] = -16'd34;
assign W_R_STAGE_LUT[1962] = -16'd254;
assign W_I_STAGE_LUT[1962] = -16'd34;
assign W_R_STAGE_LUT[1963] = -16'd254;
assign W_I_STAGE_LUT[1963] = -16'd33;
assign W_R_STAGE_LUT[1964] = -16'd254;
assign W_I_STAGE_LUT[1964] = -16'd33;
assign W_R_STAGE_LUT[1965] = -16'd254;
assign W_I_STAGE_LUT[1965] = -16'd33;
assign W_R_STAGE_LUT[1966] = -16'd254;
assign W_I_STAGE_LUT[1966] = -16'd32;
assign W_R_STAGE_LUT[1967] = -16'd254;
assign W_I_STAGE_LUT[1967] = -16'd32;
assign W_R_STAGE_LUT[1968] = -16'd254;
assign W_I_STAGE_LUT[1968] = -16'd31;
assign W_R_STAGE_LUT[1969] = -16'd254;
assign W_I_STAGE_LUT[1969] = -16'd31;
assign W_R_STAGE_LUT[1970] = -16'd254;
assign W_I_STAGE_LUT[1970] = -16'd31;
assign W_R_STAGE_LUT[1971] = -16'd254;
assign W_I_STAGE_LUT[1971] = -16'd30;
assign W_R_STAGE_LUT[1972] = -16'd254;
assign W_I_STAGE_LUT[1972] = -16'd30;
assign W_R_STAGE_LUT[1973] = -16'd254;
assign W_I_STAGE_LUT[1973] = -16'd29;
assign W_R_STAGE_LUT[1974] = -16'd254;
assign W_I_STAGE_LUT[1974] = -16'd29;
assign W_R_STAGE_LUT[1975] = -16'd254;
assign W_I_STAGE_LUT[1975] = -16'd29;
assign W_R_STAGE_LUT[1976] = -16'd254;
assign W_I_STAGE_LUT[1976] = -16'd28;
assign W_R_STAGE_LUT[1977] = -16'd254;
assign W_I_STAGE_LUT[1977] = -16'd28;
assign W_R_STAGE_LUT[1978] = -16'd255;
assign W_I_STAGE_LUT[1978] = -16'd27;
assign W_R_STAGE_LUT[1979] = -16'd255;
assign W_I_STAGE_LUT[1979] = -16'd27;
assign W_R_STAGE_LUT[1980] = -16'd255;
assign W_I_STAGE_LUT[1980] = -16'd27;
assign W_R_STAGE_LUT[1981] = -16'd255;
assign W_I_STAGE_LUT[1981] = -16'd26;
assign W_R_STAGE_LUT[1982] = -16'd255;
assign W_I_STAGE_LUT[1982] = -16'd26;
assign W_R_STAGE_LUT[1983] = -16'd255;
assign W_I_STAGE_LUT[1983] = -16'd25;
assign W_R_STAGE_LUT[1984] = -16'd255;
assign W_I_STAGE_LUT[1984] = -16'd25;
assign W_R_STAGE_LUT[1985] = -16'd255;
assign W_I_STAGE_LUT[1985] = -16'd25;
assign W_R_STAGE_LUT[1986] = -16'd255;
assign W_I_STAGE_LUT[1986] = -16'd24;
assign W_R_STAGE_LUT[1987] = -16'd255;
assign W_I_STAGE_LUT[1987] = -16'd24;
assign W_R_STAGE_LUT[1988] = -16'd255;
assign W_I_STAGE_LUT[1988] = -16'd24;
assign W_R_STAGE_LUT[1989] = -16'd255;
assign W_I_STAGE_LUT[1989] = -16'd23;
assign W_R_STAGE_LUT[1990] = -16'd255;
assign W_I_STAGE_LUT[1990] = -16'd23;
assign W_R_STAGE_LUT[1991] = -16'd255;
assign W_I_STAGE_LUT[1991] = -16'd22;
assign W_R_STAGE_LUT[1992] = -16'd255;
assign W_I_STAGE_LUT[1992] = -16'd22;
assign W_R_STAGE_LUT[1993] = -16'd255;
assign W_I_STAGE_LUT[1993] = -16'd22;
assign W_R_STAGE_LUT[1994] = -16'd255;
assign W_I_STAGE_LUT[1994] = -16'd21;
assign W_R_STAGE_LUT[1995] = -16'd255;
assign W_I_STAGE_LUT[1995] = -16'd21;
assign W_R_STAGE_LUT[1996] = -16'd255;
assign W_I_STAGE_LUT[1996] = -16'd20;
assign W_R_STAGE_LUT[1997] = -16'd255;
assign W_I_STAGE_LUT[1997] = -16'd20;
assign W_R_STAGE_LUT[1998] = -16'd255;
assign W_I_STAGE_LUT[1998] = -16'd20;
assign W_R_STAGE_LUT[1999] = -16'd255;
assign W_I_STAGE_LUT[1999] = -16'd19;
assign W_R_STAGE_LUT[2000] = -16'd255;
assign W_I_STAGE_LUT[2000] = -16'd19;
assign W_R_STAGE_LUT[2001] = -16'd255;
assign W_I_STAGE_LUT[2001] = -16'd18;
assign W_R_STAGE_LUT[2002] = -16'd255;
assign W_I_STAGE_LUT[2002] = -16'd18;
assign W_R_STAGE_LUT[2003] = -16'd255;
assign W_I_STAGE_LUT[2003] = -16'd18;
assign W_R_STAGE_LUT[2004] = -16'd255;
assign W_I_STAGE_LUT[2004] = -16'd17;
assign W_R_STAGE_LUT[2005] = -16'd255;
assign W_I_STAGE_LUT[2005] = -16'd17;
assign W_R_STAGE_LUT[2006] = -16'd255;
assign W_I_STAGE_LUT[2006] = -16'd16;
assign W_R_STAGE_LUT[2007] = -16'd255;
assign W_I_STAGE_LUT[2007] = -16'd16;
assign W_R_STAGE_LUT[2008] = -16'd256;
assign W_I_STAGE_LUT[2008] = -16'd16;
assign W_R_STAGE_LUT[2009] = -16'd256;
assign W_I_STAGE_LUT[2009] = -16'd15;
assign W_R_STAGE_LUT[2010] = -16'd256;
assign W_I_STAGE_LUT[2010] = -16'd15;
assign W_R_STAGE_LUT[2011] = -16'd256;
assign W_I_STAGE_LUT[2011] = -16'd15;
assign W_R_STAGE_LUT[2012] = -16'd256;
assign W_I_STAGE_LUT[2012] = -16'd14;
assign W_R_STAGE_LUT[2013] = -16'd256;
assign W_I_STAGE_LUT[2013] = -16'd14;
assign W_R_STAGE_LUT[2014] = -16'd256;
assign W_I_STAGE_LUT[2014] = -16'd13;
assign W_R_STAGE_LUT[2015] = -16'd256;
assign W_I_STAGE_LUT[2015] = -16'd13;
assign W_R_STAGE_LUT[2016] = -16'd256;
assign W_I_STAGE_LUT[2016] = -16'd13;
assign W_R_STAGE_LUT[2017] = -16'd256;
assign W_I_STAGE_LUT[2017] = -16'd12;
assign W_R_STAGE_LUT[2018] = -16'd256;
assign W_I_STAGE_LUT[2018] = -16'd12;
assign W_R_STAGE_LUT[2019] = -16'd256;
assign W_I_STAGE_LUT[2019] = -16'd11;
assign W_R_STAGE_LUT[2020] = -16'd256;
assign W_I_STAGE_LUT[2020] = -16'd11;
assign W_R_STAGE_LUT[2021] = -16'd256;
assign W_I_STAGE_LUT[2021] = -16'd11;
assign W_R_STAGE_LUT[2022] = -16'd256;
assign W_I_STAGE_LUT[2022] = -16'd10;
assign W_R_STAGE_LUT[2023] = -16'd256;
assign W_I_STAGE_LUT[2023] = -16'd10;
assign W_R_STAGE_LUT[2024] = -16'd256;
assign W_I_STAGE_LUT[2024] = -16'd9;
assign W_R_STAGE_LUT[2025] = -16'd256;
assign W_I_STAGE_LUT[2025] = -16'd9;
assign W_R_STAGE_LUT[2026] = -16'd256;
assign W_I_STAGE_LUT[2026] = -16'd9;
assign W_R_STAGE_LUT[2027] = -16'd256;
assign W_I_STAGE_LUT[2027] = -16'd8;
assign W_R_STAGE_LUT[2028] = -16'd256;
assign W_I_STAGE_LUT[2028] = -16'd8;
assign W_R_STAGE_LUT[2029] = -16'd256;
assign W_I_STAGE_LUT[2029] = -16'd7;
assign W_R_STAGE_LUT[2030] = -16'd256;
assign W_I_STAGE_LUT[2030] = -16'd7;
assign W_R_STAGE_LUT[2031] = -16'd256;
assign W_I_STAGE_LUT[2031] = -16'd7;
assign W_R_STAGE_LUT[2032] = -16'd256;
assign W_I_STAGE_LUT[2032] = -16'd6;
assign W_R_STAGE_LUT[2033] = -16'd256;
assign W_I_STAGE_LUT[2033] = -16'd6;
assign W_R_STAGE_LUT[2034] = -16'd256;
assign W_I_STAGE_LUT[2034] = -16'd5;
assign W_R_STAGE_LUT[2035] = -16'd256;
assign W_I_STAGE_LUT[2035] = -16'd5;
assign W_R_STAGE_LUT[2036] = -16'd256;
assign W_I_STAGE_LUT[2036] = -16'd5;
assign W_R_STAGE_LUT[2037] = -16'd256;
assign W_I_STAGE_LUT[2037] = -16'd4;
assign W_R_STAGE_LUT[2038] = -16'd256;
assign W_I_STAGE_LUT[2038] = -16'd4;
assign W_R_STAGE_LUT[2039] = -16'd256;
assign W_I_STAGE_LUT[2039] = -16'd4;
assign W_R_STAGE_LUT[2040] = -16'd256;
assign W_I_STAGE_LUT[2040] = -16'd3;
assign W_R_STAGE_LUT[2041] = -16'd256;
assign W_I_STAGE_LUT[2041] = -16'd3;
assign W_R_STAGE_LUT[2042] = -16'd256;
assign W_I_STAGE_LUT[2042] = -16'd2;
assign W_R_STAGE_LUT[2043] = -16'd256;
assign W_I_STAGE_LUT[2043] = -16'd2;
assign W_R_STAGE_LUT[2044] = -16'd256;
assign W_I_STAGE_LUT[2044] = -16'd2;
assign W_R_STAGE_LUT[2045] = -16'd256;
assign W_I_STAGE_LUT[2045] = -16'd1;
assign W_R_STAGE_LUT[2046] = -16'd256;
assign W_I_STAGE_LUT[2046] = -16'd1;
assign W_R_STAGE_LUT[2047] = -16'd256;
assign W_I_STAGE_LUT[2047] = 16'd0;
