// In the delay commutator, for each stage, delay by N/k samples where k ranges from 4 to N in powers of two.