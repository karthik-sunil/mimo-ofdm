module fft_rad2();

// N = 8 Point DIF FFT

// Using a pipelined design from lecture
// Log2(N) = 3 butterfly stages
// Each stage takes N/2 cycles

// Stage 1
// Butterfly 1
// Delay Commutator - Delay and rearrage stage output

// Stage 2
// Butterfly 2
// Delay Commutator - Delay and rearrage stage output

// Stage 3
// Butterfly 3
// Delay Commutator - Delay and rearrage stage output

endmodule