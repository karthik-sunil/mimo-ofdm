assign W_R_STAGE_LUT[0] =  16'd256; assign W_I_STAGE_LUT[0] =   16'd0;
assign W_R_STAGE_LUT[1] =  16'd237; assign W_I_STAGE_LUT[1] =  -16'd98;
assign W_R_STAGE_LUT[2] =  16'd181; assign W_I_STAGE_LUT[2] = -16'd181;
assign W_R_STAGE_LUT[3] =   16'd98; assign W_I_STAGE_LUT[3] = -16'd237;
assign W_R_STAGE_LUT[4] =    16'd0; assign W_I_STAGE_LUT[4] = -16'd256;
assign W_R_STAGE_LUT[5] =  -16'd98; assign W_I_STAGE_LUT[5] = -16'd237;
assign W_R_STAGE_LUT[6] = -16'd181; assign W_I_STAGE_LUT[6] = -16'd181;
assign W_R_STAGE_LUT[7] = -16'd237; assign W_I_STAGE_LUT[7] =  -16'd98;