assign W_R_STAGE_LUT[0]  =  16'd256; assign W_I_STAGE_LUT[0]  =    16'd0;
assign W_R_STAGE_LUT[1]  =  16'd256; assign W_I_STAGE_LUT[1]  =  -16'd13;
assign W_R_STAGE_LUT[2]  =  16'd255; assign W_I_STAGE_LUT[2]  =  -16'd25;
assign W_R_STAGE_LUT[3]  =  16'd253; assign W_I_STAGE_LUT[3]  =  -16'd38;
assign W_R_STAGE_LUT[4]  =  16'd251; assign W_I_STAGE_LUT[4]  =  -16'd50;
assign W_R_STAGE_LUT[5]  =  16'd248; assign W_I_STAGE_LUT[5]  =  -16'd62;
assign W_R_STAGE_LUT[6]  =  16'd245; assign W_I_STAGE_LUT[6]  =  -16'd74;
assign W_R_STAGE_LUT[7]  =  16'd241; assign W_I_STAGE_LUT[7]  =  -16'd86;
assign W_R_STAGE_LUT[8]  =  16'd237; assign W_I_STAGE_LUT[8]  =  -16'd98;
assign W_R_STAGE_LUT[9]  =  16'd231; assign W_I_STAGE_LUT[9]  = -16'd109;
assign W_R_STAGE_LUT[10] =  16'd226; assign W_I_STAGE_LUT[10] = -16'd121;
assign W_R_STAGE_LUT[11] =  16'd220; assign W_I_STAGE_LUT[11] = -16'd132;
assign W_R_STAGE_LUT[12] =  16'd213; assign W_I_STAGE_LUT[12] = -16'd142;
assign W_R_STAGE_LUT[13] =  16'd206; assign W_I_STAGE_LUT[13] = -16'd152;
assign W_R_STAGE_LUT[14] =  16'd198; assign W_I_STAGE_LUT[14] = -16'd162;
assign W_R_STAGE_LUT[15] =  16'd190; assign W_I_STAGE_LUT[15] = -16'd172;
assign W_R_STAGE_LUT[16] =  16'd181; assign W_I_STAGE_LUT[16] = -16'd181;
assign W_R_STAGE_LUT[17] =  16'd172; assign W_I_STAGE_LUT[17] = -16'd190;
assign W_R_STAGE_LUT[18] =  16'd162; assign W_I_STAGE_LUT[18] = -16'd198;
assign W_R_STAGE_LUT[19] =  16'd152; assign W_I_STAGE_LUT[19] = -16'd206;
assign W_R_STAGE_LUT[20] =  16'd142; assign W_I_STAGE_LUT[20] = -16'd213;
assign W_R_STAGE_LUT[21] =  16'd132; assign W_I_STAGE_LUT[21] = -16'd220;
assign W_R_STAGE_LUT[22] =  16'd121; assign W_I_STAGE_LUT[22] = -16'd226;
assign W_R_STAGE_LUT[23] =  16'd109; assign W_I_STAGE_LUT[23] = -16'd231;
assign W_R_STAGE_LUT[24] =   16'd98; assign W_I_STAGE_LUT[24] = -16'd237;
assign W_R_STAGE_LUT[25] =   16'd86; assign W_I_STAGE_LUT[25] = -16'd241;
assign W_R_STAGE_LUT[26] =   16'd74; assign W_I_STAGE_LUT[26] = -16'd245;
assign W_R_STAGE_LUT[27] =   16'd62; assign W_I_STAGE_LUT[27] = -16'd248;
assign W_R_STAGE_LUT[28] =   16'd50; assign W_I_STAGE_LUT[28] = -16'd251;
assign W_R_STAGE_LUT[29] =   16'd38; assign W_I_STAGE_LUT[29] = -16'd253;
assign W_R_STAGE_LUT[30] =   16'd25; assign W_I_STAGE_LUT[30] = -16'd255;
assign W_R_STAGE_LUT[31] =   16'd13; assign W_I_STAGE_LUT[31] = -16'd256;
assign W_R_STAGE_LUT[32] =    16'd0; assign W_I_STAGE_LUT[32] = -16'd256;
assign W_R_STAGE_LUT[33] =  -16'd13; assign W_I_STAGE_LUT[33] = -16'd256;
assign W_R_STAGE_LUT[34] =  -16'd25; assign W_I_STAGE_LUT[34] = -16'd255;
assign W_R_STAGE_LUT[35] =  -16'd38; assign W_I_STAGE_LUT[35] = -16'd253;
assign W_R_STAGE_LUT[36] =  -16'd50; assign W_I_STAGE_LUT[36] = -16'd251;
assign W_R_STAGE_LUT[37] =  -16'd62; assign W_I_STAGE_LUT[37] = -16'd248;
assign W_R_STAGE_LUT[38] =  -16'd74; assign W_I_STAGE_LUT[38] = -16'd245;
assign W_R_STAGE_LUT[39] =  -16'd86; assign W_I_STAGE_LUT[39] = -16'd241;
assign W_R_STAGE_LUT[40] =  -16'd98; assign W_I_STAGE_LUT[40] = -16'd237;
assign W_R_STAGE_LUT[41] = -16'd109; assign W_I_STAGE_LUT[41] = -16'd231;
assign W_R_STAGE_LUT[42] = -16'd121; assign W_I_STAGE_LUT[42] = -16'd226;
assign W_R_STAGE_LUT[43] = -16'd132; assign W_I_STAGE_LUT[43] = -16'd220;
assign W_R_STAGE_LUT[44] = -16'd142; assign W_I_STAGE_LUT[44] = -16'd213;
assign W_R_STAGE_LUT[45] = -16'd152; assign W_I_STAGE_LUT[45] = -16'd206;
assign W_R_STAGE_LUT[46] = -16'd162; assign W_I_STAGE_LUT[46] = -16'd198;
assign W_R_STAGE_LUT[47] = -16'd172; assign W_I_STAGE_LUT[47] = -16'd190;
assign W_R_STAGE_LUT[48] = -16'd181; assign W_I_STAGE_LUT[48] = -16'd181;
assign W_R_STAGE_LUT[49] = -16'd190; assign W_I_STAGE_LUT[49] = -16'd172;
assign W_R_STAGE_LUT[50] = -16'd198; assign W_I_STAGE_LUT[50] = -16'd162;
assign W_R_STAGE_LUT[51] = -16'd206; assign W_I_STAGE_LUT[51] = -16'd152;
assign W_R_STAGE_LUT[52] = -16'd213; assign W_I_STAGE_LUT[52] = -16'd142;
assign W_R_STAGE_LUT[53] = -16'd220; assign W_I_STAGE_LUT[53] = -16'd132;
assign W_R_STAGE_LUT[54] = -16'd226; assign W_I_STAGE_LUT[54] = -16'd121;
assign W_R_STAGE_LUT[55] = -16'd231; assign W_I_STAGE_LUT[55] = -16'd109;
assign W_R_STAGE_LUT[56] = -16'd237; assign W_I_STAGE_LUT[56] =  -16'd98;
assign W_R_STAGE_LUT[57] = -16'd241; assign W_I_STAGE_LUT[57] =  -16'd86;
assign W_R_STAGE_LUT[58] = -16'd245; assign W_I_STAGE_LUT[58] =  -16'd74;
assign W_R_STAGE_LUT[59] = -16'd248; assign W_I_STAGE_LUT[59] =  -16'd62;
assign W_R_STAGE_LUT[60] = -16'd251; assign W_I_STAGE_LUT[60] =  -16'd50;
assign W_R_STAGE_LUT[61] = -16'd253; assign W_I_STAGE_LUT[61] =  -16'd38;
assign W_R_STAGE_LUT[62] = -16'd255; assign W_I_STAGE_LUT[62] =  -16'd25;
assign W_R_STAGE_LUT[63] = -16'd256; assign W_I_STAGE_LUT[63] =  -16'd13;
