assign W_R_STAGE_LUT[0] =  256;      assign W_I_STAGE_LUT[0] =    0;
assign W_R_STAGE_LUT[1] =  181;      assign W_I_STAGE_LUT[1] = -181;
assign W_R_STAGE_LUT[2] =    0;      assign W_I_STAGE_LUT[2] = -256;
assign W_R_STAGE_LUT[3] = -181;      assign W_I_STAGE_LUT[3] = -181; 