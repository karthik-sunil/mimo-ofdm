assign W_R_STAGE_LUT[0] = 16'd256;
assign W_I_STAGE_LUT[0] = 16'd0;
assign W_R_STAGE_LUT[1] = 16'd256;
assign W_I_STAGE_LUT[1] = -16'd1;
assign W_R_STAGE_LUT[2] = 16'd256;
assign W_I_STAGE_LUT[2] = -16'd2;
assign W_R_STAGE_LUT[3] = 16'd256;
assign W_I_STAGE_LUT[3] = -16'd2;
assign W_R_STAGE_LUT[4] = 16'd256;
assign W_I_STAGE_LUT[4] = -16'd3;
assign W_R_STAGE_LUT[5] = 16'd256;
assign W_I_STAGE_LUT[5] = -16'd4;
assign W_R_STAGE_LUT[6] = 16'd256;
assign W_I_STAGE_LUT[6] = -16'd5;
assign W_R_STAGE_LUT[7] = 16'd256;
assign W_I_STAGE_LUT[7] = -16'd5;
assign W_R_STAGE_LUT[8] = 16'd256;
assign W_I_STAGE_LUT[8] = -16'd6;
assign W_R_STAGE_LUT[9] = 16'd256;
assign W_I_STAGE_LUT[9] = -16'd7;
assign W_R_STAGE_LUT[10] = 16'd256;
assign W_I_STAGE_LUT[10] = -16'd8;
assign W_R_STAGE_LUT[11] = 16'd256;
assign W_I_STAGE_LUT[11] = -16'd9;
assign W_R_STAGE_LUT[12] = 16'd256;
assign W_I_STAGE_LUT[12] = -16'd9;
assign W_R_STAGE_LUT[13] = 16'd256;
assign W_I_STAGE_LUT[13] = -16'd10;
assign W_R_STAGE_LUT[14] = 16'd256;
assign W_I_STAGE_LUT[14] = -16'd11;
assign W_R_STAGE_LUT[15] = 16'd256;
assign W_I_STAGE_LUT[15] = -16'd12;
assign W_R_STAGE_LUT[16] = 16'd256;
assign W_I_STAGE_LUT[16] = -16'd13;
assign W_R_STAGE_LUT[17] = 16'd256;
assign W_I_STAGE_LUT[17] = -16'd13;
assign W_R_STAGE_LUT[18] = 16'd256;
assign W_I_STAGE_LUT[18] = -16'd14;
assign W_R_STAGE_LUT[19] = 16'd256;
assign W_I_STAGE_LUT[19] = -16'd15;
assign W_R_STAGE_LUT[20] = 16'd256;
assign W_I_STAGE_LUT[20] = -16'd16;
assign W_R_STAGE_LUT[21] = 16'd255;
assign W_I_STAGE_LUT[21] = -16'd16;
assign W_R_STAGE_LUT[22] = 16'd255;
assign W_I_STAGE_LUT[22] = -16'd17;
assign W_R_STAGE_LUT[23] = 16'd255;
assign W_I_STAGE_LUT[23] = -16'd18;
assign W_R_STAGE_LUT[24] = 16'd255;
assign W_I_STAGE_LUT[24] = -16'd19;
assign W_R_STAGE_LUT[25] = 16'd255;
assign W_I_STAGE_LUT[25] = -16'd20;
assign W_R_STAGE_LUT[26] = 16'd255;
assign W_I_STAGE_LUT[26] = -16'd20;
assign W_R_STAGE_LUT[27] = 16'd255;
assign W_I_STAGE_LUT[27] = -16'd21;
assign W_R_STAGE_LUT[28] = 16'd255;
assign W_I_STAGE_LUT[28] = -16'd22;
assign W_R_STAGE_LUT[29] = 16'd255;
assign W_I_STAGE_LUT[29] = -16'd23;
assign W_R_STAGE_LUT[30] = 16'd255;
assign W_I_STAGE_LUT[30] = -16'd24;
assign W_R_STAGE_LUT[31] = 16'd255;
assign W_I_STAGE_LUT[31] = -16'd24;
assign W_R_STAGE_LUT[32] = 16'd255;
assign W_I_STAGE_LUT[32] = -16'd25;
assign W_R_STAGE_LUT[33] = 16'd255;
assign W_I_STAGE_LUT[33] = -16'd26;
assign W_R_STAGE_LUT[34] = 16'd255;
assign W_I_STAGE_LUT[34] = -16'd27;
assign W_R_STAGE_LUT[35] = 16'd255;
assign W_I_STAGE_LUT[35] = -16'd27;
assign W_R_STAGE_LUT[36] = 16'd254;
assign W_I_STAGE_LUT[36] = -16'd28;
assign W_R_STAGE_LUT[37] = 16'd254;
assign W_I_STAGE_LUT[37] = -16'd29;
assign W_R_STAGE_LUT[38] = 16'd254;
assign W_I_STAGE_LUT[38] = -16'd30;
assign W_R_STAGE_LUT[39] = 16'd254;
assign W_I_STAGE_LUT[39] = -16'd31;
assign W_R_STAGE_LUT[40] = 16'd254;
assign W_I_STAGE_LUT[40] = -16'd31;
assign W_R_STAGE_LUT[41] = 16'd254;
assign W_I_STAGE_LUT[41] = -16'd32;
assign W_R_STAGE_LUT[42] = 16'd254;
assign W_I_STAGE_LUT[42] = -16'd33;
assign W_R_STAGE_LUT[43] = 16'd254;
assign W_I_STAGE_LUT[43] = -16'd34;
assign W_R_STAGE_LUT[44] = 16'd254;
assign W_I_STAGE_LUT[44] = -16'd34;
assign W_R_STAGE_LUT[45] = 16'd254;
assign W_I_STAGE_LUT[45] = -16'd35;
assign W_R_STAGE_LUT[46] = 16'd253;
assign W_I_STAGE_LUT[46] = -16'd36;
assign W_R_STAGE_LUT[47] = 16'd253;
assign W_I_STAGE_LUT[47] = -16'd37;
assign W_R_STAGE_LUT[48] = 16'd253;
assign W_I_STAGE_LUT[48] = -16'd38;
assign W_R_STAGE_LUT[49] = 16'd253;
assign W_I_STAGE_LUT[49] = -16'd38;
assign W_R_STAGE_LUT[50] = 16'd253;
assign W_I_STAGE_LUT[50] = -16'd39;
assign W_R_STAGE_LUT[51] = 16'd253;
assign W_I_STAGE_LUT[51] = -16'd40;
assign W_R_STAGE_LUT[52] = 16'd253;
assign W_I_STAGE_LUT[52] = -16'd41;
assign W_R_STAGE_LUT[53] = 16'd253;
assign W_I_STAGE_LUT[53] = -16'd41;
assign W_R_STAGE_LUT[54] = 16'd252;
assign W_I_STAGE_LUT[54] = -16'd42;
assign W_R_STAGE_LUT[55] = 16'd252;
assign W_I_STAGE_LUT[55] = -16'd43;
assign W_R_STAGE_LUT[56] = 16'd252;
assign W_I_STAGE_LUT[56] = -16'd44;
assign W_R_STAGE_LUT[57] = 16'd252;
assign W_I_STAGE_LUT[57] = -16'd45;
assign W_R_STAGE_LUT[58] = 16'd252;
assign W_I_STAGE_LUT[58] = -16'd45;
assign W_R_STAGE_LUT[59] = 16'd252;
assign W_I_STAGE_LUT[59] = -16'd46;
assign W_R_STAGE_LUT[60] = 16'd252;
assign W_I_STAGE_LUT[60] = -16'd47;
assign W_R_STAGE_LUT[61] = 16'd252;
assign W_I_STAGE_LUT[61] = -16'd48;
assign W_R_STAGE_LUT[62] = 16'd251;
assign W_I_STAGE_LUT[62] = -16'd48;
assign W_R_STAGE_LUT[63] = 16'd251;
assign W_I_STAGE_LUT[63] = -16'd49;
assign W_R_STAGE_LUT[64] = 16'd251;
assign W_I_STAGE_LUT[64] = -16'd50;
assign W_R_STAGE_LUT[65] = 16'd251;
assign W_I_STAGE_LUT[65] = -16'd51;
assign W_R_STAGE_LUT[66] = 16'd251;
assign W_I_STAGE_LUT[66] = -16'd51;
assign W_R_STAGE_LUT[67] = 16'd251;
assign W_I_STAGE_LUT[67] = -16'd52;
assign W_R_STAGE_LUT[68] = 16'd250;
assign W_I_STAGE_LUT[68] = -16'd53;
assign W_R_STAGE_LUT[69] = 16'd250;
assign W_I_STAGE_LUT[69] = -16'd54;
assign W_R_STAGE_LUT[70] = 16'd250;
assign W_I_STAGE_LUT[70] = -16'd55;
assign W_R_STAGE_LUT[71] = 16'd250;
assign W_I_STAGE_LUT[71] = -16'd55;
assign W_R_STAGE_LUT[72] = 16'd250;
assign W_I_STAGE_LUT[72] = -16'd56;
assign W_R_STAGE_LUT[73] = 16'd250;
assign W_I_STAGE_LUT[73] = -16'd57;
assign W_R_STAGE_LUT[74] = 16'd249;
assign W_I_STAGE_LUT[74] = -16'd58;
assign W_R_STAGE_LUT[75] = 16'd249;
assign W_I_STAGE_LUT[75] = -16'd58;
assign W_R_STAGE_LUT[76] = 16'd249;
assign W_I_STAGE_LUT[76] = -16'd59;
assign W_R_STAGE_LUT[77] = 16'd249;
assign W_I_STAGE_LUT[77] = -16'd60;
assign W_R_STAGE_LUT[78] = 16'd249;
assign W_I_STAGE_LUT[78] = -16'd61;
assign W_R_STAGE_LUT[79] = 16'd249;
assign W_I_STAGE_LUT[79] = -16'd61;
assign W_R_STAGE_LUT[80] = 16'd248;
assign W_I_STAGE_LUT[80] = -16'd62;
assign W_R_STAGE_LUT[81] = 16'd248;
assign W_I_STAGE_LUT[81] = -16'd63;
assign W_R_STAGE_LUT[82] = 16'd248;
assign W_I_STAGE_LUT[82] = -16'd64;
assign W_R_STAGE_LUT[83] = 16'd248;
assign W_I_STAGE_LUT[83] = -16'd64;
assign W_R_STAGE_LUT[84] = 16'd248;
assign W_I_STAGE_LUT[84] = -16'd65;
assign W_R_STAGE_LUT[85] = 16'd247;
assign W_I_STAGE_LUT[85] = -16'd66;
assign W_R_STAGE_LUT[86] = 16'd247;
assign W_I_STAGE_LUT[86] = -16'd67;
assign W_R_STAGE_LUT[87] = 16'd247;
assign W_I_STAGE_LUT[87] = -16'd68;
assign W_R_STAGE_LUT[88] = 16'd247;
assign W_I_STAGE_LUT[88] = -16'd68;
assign W_R_STAGE_LUT[89] = 16'd247;
assign W_I_STAGE_LUT[89] = -16'd69;
assign W_R_STAGE_LUT[90] = 16'd246;
assign W_I_STAGE_LUT[90] = -16'd70;
assign W_R_STAGE_LUT[91] = 16'd246;
assign W_I_STAGE_LUT[91] = -16'd71;
assign W_R_STAGE_LUT[92] = 16'd246;
assign W_I_STAGE_LUT[92] = -16'd71;
assign W_R_STAGE_LUT[93] = 16'd246;
assign W_I_STAGE_LUT[93] = -16'd72;
assign W_R_STAGE_LUT[94] = 16'd245;
assign W_I_STAGE_LUT[94] = -16'd73;
assign W_R_STAGE_LUT[95] = 16'd245;
assign W_I_STAGE_LUT[95] = -16'd74;
assign W_R_STAGE_LUT[96] = 16'd245;
assign W_I_STAGE_LUT[96] = -16'd74;
assign W_R_STAGE_LUT[97] = 16'd245;
assign W_I_STAGE_LUT[97] = -16'd75;
assign W_R_STAGE_LUT[98] = 16'd245;
assign W_I_STAGE_LUT[98] = -16'd76;
assign W_R_STAGE_LUT[99] = 16'd244;
assign W_I_STAGE_LUT[99] = -16'd77;
assign W_R_STAGE_LUT[100] = 16'd244;
assign W_I_STAGE_LUT[100] = -16'd77;
assign W_R_STAGE_LUT[101] = 16'd244;
assign W_I_STAGE_LUT[101] = -16'd78;
assign W_R_STAGE_LUT[102] = 16'd244;
assign W_I_STAGE_LUT[102] = -16'd79;
assign W_R_STAGE_LUT[103] = 16'd243;
assign W_I_STAGE_LUT[103] = -16'd80;
assign W_R_STAGE_LUT[104] = 16'd243;
assign W_I_STAGE_LUT[104] = -16'd80;
assign W_R_STAGE_LUT[105] = 16'd243;
assign W_I_STAGE_LUT[105] = -16'd81;
assign W_R_STAGE_LUT[106] = 16'd243;
assign W_I_STAGE_LUT[106] = -16'd82;
assign W_R_STAGE_LUT[107] = 16'd242;
assign W_I_STAGE_LUT[107] = -16'd83;
assign W_R_STAGE_LUT[108] = 16'd242;
assign W_I_STAGE_LUT[108] = -16'd83;
assign W_R_STAGE_LUT[109] = 16'd242;
assign W_I_STAGE_LUT[109] = -16'd84;
assign W_R_STAGE_LUT[110] = 16'd242;
assign W_I_STAGE_LUT[110] = -16'd85;
assign W_R_STAGE_LUT[111] = 16'd241;
assign W_I_STAGE_LUT[111] = -16'd86;
assign W_R_STAGE_LUT[112] = 16'd241;
assign W_I_STAGE_LUT[112] = -16'd86;
assign W_R_STAGE_LUT[113] = 16'd241;
assign W_I_STAGE_LUT[113] = -16'd87;
assign W_R_STAGE_LUT[114] = 16'd241;
assign W_I_STAGE_LUT[114] = -16'd88;
assign W_R_STAGE_LUT[115] = 16'd240;
assign W_I_STAGE_LUT[115] = -16'd88;
assign W_R_STAGE_LUT[116] = 16'd240;
assign W_I_STAGE_LUT[116] = -16'd89;
assign W_R_STAGE_LUT[117] = 16'd240;
assign W_I_STAGE_LUT[117] = -16'd90;
assign W_R_STAGE_LUT[118] = 16'd239;
assign W_I_STAGE_LUT[118] = -16'd91;
assign W_R_STAGE_LUT[119] = 16'd239;
assign W_I_STAGE_LUT[119] = -16'd91;
assign W_R_STAGE_LUT[120] = 16'd239;
assign W_I_STAGE_LUT[120] = -16'd92;
assign W_R_STAGE_LUT[121] = 16'd239;
assign W_I_STAGE_LUT[121] = -16'd93;
assign W_R_STAGE_LUT[122] = 16'd238;
assign W_I_STAGE_LUT[122] = -16'd94;
assign W_R_STAGE_LUT[123] = 16'd238;
assign W_I_STAGE_LUT[123] = -16'd94;
assign W_R_STAGE_LUT[124] = 16'd238;
assign W_I_STAGE_LUT[124] = -16'd95;
assign W_R_STAGE_LUT[125] = 16'd237;
assign W_I_STAGE_LUT[125] = -16'd96;
assign W_R_STAGE_LUT[126] = 16'd237;
assign W_I_STAGE_LUT[126] = -16'd97;
assign W_R_STAGE_LUT[127] = 16'd237;
assign W_I_STAGE_LUT[127] = -16'd97;
assign W_R_STAGE_LUT[128] = 16'd237;
assign W_I_STAGE_LUT[128] = -16'd98;
assign W_R_STAGE_LUT[129] = 16'd236;
assign W_I_STAGE_LUT[129] = -16'd99;
assign W_R_STAGE_LUT[130] = 16'd236;
assign W_I_STAGE_LUT[130] = -16'd99;
assign W_R_STAGE_LUT[131] = 16'd236;
assign W_I_STAGE_LUT[131] = -16'd100;
assign W_R_STAGE_LUT[132] = 16'd235;
assign W_I_STAGE_LUT[132] = -16'd101;
assign W_R_STAGE_LUT[133] = 16'd235;
assign W_I_STAGE_LUT[133] = -16'd102;
assign W_R_STAGE_LUT[134] = 16'd235;
assign W_I_STAGE_LUT[134] = -16'd102;
assign W_R_STAGE_LUT[135] = 16'd234;
assign W_I_STAGE_LUT[135] = -16'd103;
assign W_R_STAGE_LUT[136] = 16'd234;
assign W_I_STAGE_LUT[136] = -16'd104;
assign W_R_STAGE_LUT[137] = 16'd234;
assign W_I_STAGE_LUT[137] = -16'd104;
assign W_R_STAGE_LUT[138] = 16'd233;
assign W_I_STAGE_LUT[138] = -16'd105;
assign W_R_STAGE_LUT[139] = 16'd233;
assign W_I_STAGE_LUT[139] = -16'd106;
assign W_R_STAGE_LUT[140] = 16'd233;
assign W_I_STAGE_LUT[140] = -16'd107;
assign W_R_STAGE_LUT[141] = 16'd232;
assign W_I_STAGE_LUT[141] = -16'd107;
assign W_R_STAGE_LUT[142] = 16'd232;
assign W_I_STAGE_LUT[142] = -16'd108;
assign W_R_STAGE_LUT[143] = 16'd232;
assign W_I_STAGE_LUT[143] = -16'd109;
assign W_R_STAGE_LUT[144] = 16'd231;
assign W_I_STAGE_LUT[144] = -16'd109;
assign W_R_STAGE_LUT[145] = 16'd231;
assign W_I_STAGE_LUT[145] = -16'd110;
assign W_R_STAGE_LUT[146] = 16'd231;
assign W_I_STAGE_LUT[146] = -16'd111;
assign W_R_STAGE_LUT[147] = 16'd230;
assign W_I_STAGE_LUT[147] = -16'd112;
assign W_R_STAGE_LUT[148] = 16'd230;
assign W_I_STAGE_LUT[148] = -16'd112;
assign W_R_STAGE_LUT[149] = 16'd230;
assign W_I_STAGE_LUT[149] = -16'd113;
assign W_R_STAGE_LUT[150] = 16'd229;
assign W_I_STAGE_LUT[150] = -16'd114;
assign W_R_STAGE_LUT[151] = 16'd229;
assign W_I_STAGE_LUT[151] = -16'd114;
assign W_R_STAGE_LUT[152] = 16'd229;
assign W_I_STAGE_LUT[152] = -16'd115;
assign W_R_STAGE_LUT[153] = 16'd228;
assign W_I_STAGE_LUT[153] = -16'd116;
assign W_R_STAGE_LUT[154] = 16'd228;
assign W_I_STAGE_LUT[154] = -16'd117;
assign W_R_STAGE_LUT[155] = 16'd228;
assign W_I_STAGE_LUT[155] = -16'd117;
assign W_R_STAGE_LUT[156] = 16'd227;
assign W_I_STAGE_LUT[156] = -16'd118;
assign W_R_STAGE_LUT[157] = 16'd227;
assign W_I_STAGE_LUT[157] = -16'd119;
assign W_R_STAGE_LUT[158] = 16'd227;
assign W_I_STAGE_LUT[158] = -16'd119;
assign W_R_STAGE_LUT[159] = 16'd226;
assign W_I_STAGE_LUT[159] = -16'd120;
assign W_R_STAGE_LUT[160] = 16'd226;
assign W_I_STAGE_LUT[160] = -16'd121;
assign W_R_STAGE_LUT[161] = 16'd225;
assign W_I_STAGE_LUT[161] = -16'd121;
assign W_R_STAGE_LUT[162] = 16'd225;
assign W_I_STAGE_LUT[162] = -16'd122;
assign W_R_STAGE_LUT[163] = 16'd225;
assign W_I_STAGE_LUT[163] = -16'd123;
assign W_R_STAGE_LUT[164] = 16'd224;
assign W_I_STAGE_LUT[164] = -16'd123;
assign W_R_STAGE_LUT[165] = 16'd224;
assign W_I_STAGE_LUT[165] = -16'd124;
assign W_R_STAGE_LUT[166] = 16'd224;
assign W_I_STAGE_LUT[166] = -16'd125;
assign W_R_STAGE_LUT[167] = 16'd223;
assign W_I_STAGE_LUT[167] = -16'd125;
assign W_R_STAGE_LUT[168] = 16'd223;
assign W_I_STAGE_LUT[168] = -16'd126;
assign W_R_STAGE_LUT[169] = 16'd222;
assign W_I_STAGE_LUT[169] = -16'd127;
assign W_R_STAGE_LUT[170] = 16'd222;
assign W_I_STAGE_LUT[170] = -16'd128;
assign W_R_STAGE_LUT[171] = 16'd222;
assign W_I_STAGE_LUT[171] = -16'd128;
assign W_R_STAGE_LUT[172] = 16'd221;
assign W_I_STAGE_LUT[172] = -16'd129;
assign W_R_STAGE_LUT[173] = 16'd221;
assign W_I_STAGE_LUT[173] = -16'd130;
assign W_R_STAGE_LUT[174] = 16'd220;
assign W_I_STAGE_LUT[174] = -16'd130;
assign W_R_STAGE_LUT[175] = 16'd220;
assign W_I_STAGE_LUT[175] = -16'd131;
assign W_R_STAGE_LUT[176] = 16'd220;
assign W_I_STAGE_LUT[176] = -16'd132;
assign W_R_STAGE_LUT[177] = 16'd219;
assign W_I_STAGE_LUT[177] = -16'd132;
assign W_R_STAGE_LUT[178] = 16'd219;
assign W_I_STAGE_LUT[178] = -16'd133;
assign W_R_STAGE_LUT[179] = 16'd218;
assign W_I_STAGE_LUT[179] = -16'd134;
assign W_R_STAGE_LUT[180] = 16'd218;
assign W_I_STAGE_LUT[180] = -16'd134;
assign W_R_STAGE_LUT[181] = 16'd218;
assign W_I_STAGE_LUT[181] = -16'd135;
assign W_R_STAGE_LUT[182] = 16'd217;
assign W_I_STAGE_LUT[182] = -16'd136;
assign W_R_STAGE_LUT[183] = 16'd217;
assign W_I_STAGE_LUT[183] = -16'd136;
assign W_R_STAGE_LUT[184] = 16'd216;
assign W_I_STAGE_LUT[184] = -16'd137;
assign W_R_STAGE_LUT[185] = 16'd216;
assign W_I_STAGE_LUT[185] = -16'd138;
assign W_R_STAGE_LUT[186] = 16'd215;
assign W_I_STAGE_LUT[186] = -16'd138;
assign W_R_STAGE_LUT[187] = 16'd215;
assign W_I_STAGE_LUT[187] = -16'd139;
assign W_R_STAGE_LUT[188] = 16'd215;
assign W_I_STAGE_LUT[188] = -16'd140;
assign W_R_STAGE_LUT[189] = 16'd214;
assign W_I_STAGE_LUT[189] = -16'd140;
assign W_R_STAGE_LUT[190] = 16'd214;
assign W_I_STAGE_LUT[190] = -16'd141;
assign W_R_STAGE_LUT[191] = 16'd213;
assign W_I_STAGE_LUT[191] = -16'd142;
assign W_R_STAGE_LUT[192] = 16'd213;
assign W_I_STAGE_LUT[192] = -16'd142;
assign W_R_STAGE_LUT[193] = 16'd212;
assign W_I_STAGE_LUT[193] = -16'd143;
assign W_R_STAGE_LUT[194] = 16'd212;
assign W_I_STAGE_LUT[194] = -16'd144;
assign W_R_STAGE_LUT[195] = 16'd212;
assign W_I_STAGE_LUT[195] = -16'd144;
assign W_R_STAGE_LUT[196] = 16'd211;
assign W_I_STAGE_LUT[196] = -16'd145;
assign W_R_STAGE_LUT[197] = 16'd211;
assign W_I_STAGE_LUT[197] = -16'd145;
assign W_R_STAGE_LUT[198] = 16'd210;
assign W_I_STAGE_LUT[198] = -16'd146;
assign W_R_STAGE_LUT[199] = 16'd210;
assign W_I_STAGE_LUT[199] = -16'd147;
assign W_R_STAGE_LUT[200] = 16'd209;
assign W_I_STAGE_LUT[200] = -16'd147;
assign W_R_STAGE_LUT[201] = 16'd209;
assign W_I_STAGE_LUT[201] = -16'd148;
assign W_R_STAGE_LUT[202] = 16'd208;
assign W_I_STAGE_LUT[202] = -16'd149;
assign W_R_STAGE_LUT[203] = 16'd208;
assign W_I_STAGE_LUT[203] = -16'd149;
assign W_R_STAGE_LUT[204] = 16'd207;
assign W_I_STAGE_LUT[204] = -16'd150;
assign W_R_STAGE_LUT[205] = 16'd207;
assign W_I_STAGE_LUT[205] = -16'd151;
assign W_R_STAGE_LUT[206] = 16'd207;
assign W_I_STAGE_LUT[206] = -16'd151;
assign W_R_STAGE_LUT[207] = 16'd206;
assign W_I_STAGE_LUT[207] = -16'd152;
assign W_R_STAGE_LUT[208] = 16'd206;
assign W_I_STAGE_LUT[208] = -16'd152;
assign W_R_STAGE_LUT[209] = 16'd205;
assign W_I_STAGE_LUT[209] = -16'd153;
assign W_R_STAGE_LUT[210] = 16'd205;
assign W_I_STAGE_LUT[210] = -16'd154;
assign W_R_STAGE_LUT[211] = 16'd204;
assign W_I_STAGE_LUT[211] = -16'd154;
assign W_R_STAGE_LUT[212] = 16'd204;
assign W_I_STAGE_LUT[212] = -16'd155;
assign W_R_STAGE_LUT[213] = 16'd203;
assign W_I_STAGE_LUT[213] = -16'd156;
assign W_R_STAGE_LUT[214] = 16'd203;
assign W_I_STAGE_LUT[214] = -16'd156;
assign W_R_STAGE_LUT[215] = 16'd202;
assign W_I_STAGE_LUT[215] = -16'd157;
assign W_R_STAGE_LUT[216] = 16'd202;
assign W_I_STAGE_LUT[216] = -16'd157;
assign W_R_STAGE_LUT[217] = 16'd201;
assign W_I_STAGE_LUT[217] = -16'd158;
assign W_R_STAGE_LUT[218] = 16'd201;
assign W_I_STAGE_LUT[218] = -16'd159;
assign W_R_STAGE_LUT[219] = 16'd200;
assign W_I_STAGE_LUT[219] = -16'd159;
assign W_R_STAGE_LUT[220] = 16'd200;
assign W_I_STAGE_LUT[220] = -16'd160;
assign W_R_STAGE_LUT[221] = 16'd199;
assign W_I_STAGE_LUT[221] = -16'd161;
assign W_R_STAGE_LUT[222] = 16'd199;
assign W_I_STAGE_LUT[222] = -16'd161;
assign W_R_STAGE_LUT[223] = 16'd198;
assign W_I_STAGE_LUT[223] = -16'd162;
assign W_R_STAGE_LUT[224] = 16'd198;
assign W_I_STAGE_LUT[224] = -16'd162;
assign W_R_STAGE_LUT[225] = 16'd197;
assign W_I_STAGE_LUT[225] = -16'd163;
assign W_R_STAGE_LUT[226] = 16'd197;
assign W_I_STAGE_LUT[226] = -16'd164;
assign W_R_STAGE_LUT[227] = 16'd196;
assign W_I_STAGE_LUT[227] = -16'd164;
assign W_R_STAGE_LUT[228] = 16'd196;
assign W_I_STAGE_LUT[228] = -16'd165;
assign W_R_STAGE_LUT[229] = 16'd195;
assign W_I_STAGE_LUT[229] = -16'd165;
assign W_R_STAGE_LUT[230] = 16'd195;
assign W_I_STAGE_LUT[230] = -16'd166;
assign W_R_STAGE_LUT[231] = 16'd194;
assign W_I_STAGE_LUT[231] = -16'd167;
assign W_R_STAGE_LUT[232] = 16'd194;
assign W_I_STAGE_LUT[232] = -16'd167;
assign W_R_STAGE_LUT[233] = 16'd193;
assign W_I_STAGE_LUT[233] = -16'd168;
assign W_R_STAGE_LUT[234] = 16'd193;
assign W_I_STAGE_LUT[234] = -16'd168;
assign W_R_STAGE_LUT[235] = 16'd192;
assign W_I_STAGE_LUT[235] = -16'd169;
assign W_R_STAGE_LUT[236] = 16'd192;
assign W_I_STAGE_LUT[236] = -16'd170;
assign W_R_STAGE_LUT[237] = 16'd191;
assign W_I_STAGE_LUT[237] = -16'd170;
assign W_R_STAGE_LUT[238] = 16'd191;
assign W_I_STAGE_LUT[238] = -16'd171;
assign W_R_STAGE_LUT[239] = 16'd190;
assign W_I_STAGE_LUT[239] = -16'd171;
assign W_R_STAGE_LUT[240] = 16'd190;
assign W_I_STAGE_LUT[240] = -16'd172;
assign W_R_STAGE_LUT[241] = 16'd189;
assign W_I_STAGE_LUT[241] = -16'd173;
assign W_R_STAGE_LUT[242] = 16'd189;
assign W_I_STAGE_LUT[242] = -16'd173;
assign W_R_STAGE_LUT[243] = 16'd188;
assign W_I_STAGE_LUT[243] = -16'd174;
assign W_R_STAGE_LUT[244] = 16'd188;
assign W_I_STAGE_LUT[244] = -16'd174;
assign W_R_STAGE_LUT[245] = 16'd187;
assign W_I_STAGE_LUT[245] = -16'd175;
assign W_R_STAGE_LUT[246] = 16'd186;
assign W_I_STAGE_LUT[246] = -16'd175;
assign W_R_STAGE_LUT[247] = 16'd186;
assign W_I_STAGE_LUT[247] = -16'd176;
assign W_R_STAGE_LUT[248] = 16'd185;
assign W_I_STAGE_LUT[248] = -16'd177;
assign W_R_STAGE_LUT[249] = 16'd185;
assign W_I_STAGE_LUT[249] = -16'd177;
assign W_R_STAGE_LUT[250] = 16'd184;
assign W_I_STAGE_LUT[250] = -16'd178;
assign W_R_STAGE_LUT[251] = 16'd184;
assign W_I_STAGE_LUT[251] = -16'd178;
assign W_R_STAGE_LUT[252] = 16'd183;
assign W_I_STAGE_LUT[252] = -16'd179;
assign W_R_STAGE_LUT[253] = 16'd183;
assign W_I_STAGE_LUT[253] = -16'd179;
assign W_R_STAGE_LUT[254] = 16'd182;
assign W_I_STAGE_LUT[254] = -16'd180;
assign W_R_STAGE_LUT[255] = 16'd182;
assign W_I_STAGE_LUT[255] = -16'd180;
assign W_R_STAGE_LUT[256] = 16'd181;
assign W_I_STAGE_LUT[256] = -16'd181;
assign W_R_STAGE_LUT[257] = 16'd180;
assign W_I_STAGE_LUT[257] = -16'd182;
assign W_R_STAGE_LUT[258] = 16'd180;
assign W_I_STAGE_LUT[258] = -16'd182;
assign W_R_STAGE_LUT[259] = 16'd179;
assign W_I_STAGE_LUT[259] = -16'd183;
assign W_R_STAGE_LUT[260] = 16'd179;
assign W_I_STAGE_LUT[260] = -16'd183;
assign W_R_STAGE_LUT[261] = 16'd178;
assign W_I_STAGE_LUT[261] = -16'd184;
assign W_R_STAGE_LUT[262] = 16'd178;
assign W_I_STAGE_LUT[262] = -16'd184;
assign W_R_STAGE_LUT[263] = 16'd177;
assign W_I_STAGE_LUT[263] = -16'd185;
assign W_R_STAGE_LUT[264] = 16'd177;
assign W_I_STAGE_LUT[264] = -16'd185;
assign W_R_STAGE_LUT[265] = 16'd176;
assign W_I_STAGE_LUT[265] = -16'd186;
assign W_R_STAGE_LUT[266] = 16'd175;
assign W_I_STAGE_LUT[266] = -16'd186;
assign W_R_STAGE_LUT[267] = 16'd175;
assign W_I_STAGE_LUT[267] = -16'd187;
assign W_R_STAGE_LUT[268] = 16'd174;
assign W_I_STAGE_LUT[268] = -16'd188;
assign W_R_STAGE_LUT[269] = 16'd174;
assign W_I_STAGE_LUT[269] = -16'd188;
assign W_R_STAGE_LUT[270] = 16'd173;
assign W_I_STAGE_LUT[270] = -16'd189;
assign W_R_STAGE_LUT[271] = 16'd173;
assign W_I_STAGE_LUT[271] = -16'd189;
assign W_R_STAGE_LUT[272] = 16'd172;
assign W_I_STAGE_LUT[272] = -16'd190;
assign W_R_STAGE_LUT[273] = 16'd171;
assign W_I_STAGE_LUT[273] = -16'd190;
assign W_R_STAGE_LUT[274] = 16'd171;
assign W_I_STAGE_LUT[274] = -16'd191;
assign W_R_STAGE_LUT[275] = 16'd170;
assign W_I_STAGE_LUT[275] = -16'd191;
assign W_R_STAGE_LUT[276] = 16'd170;
assign W_I_STAGE_LUT[276] = -16'd192;
assign W_R_STAGE_LUT[277] = 16'd169;
assign W_I_STAGE_LUT[277] = -16'd192;
assign W_R_STAGE_LUT[278] = 16'd168;
assign W_I_STAGE_LUT[278] = -16'd193;
assign W_R_STAGE_LUT[279] = 16'd168;
assign W_I_STAGE_LUT[279] = -16'd193;
assign W_R_STAGE_LUT[280] = 16'd167;
assign W_I_STAGE_LUT[280] = -16'd194;
assign W_R_STAGE_LUT[281] = 16'd167;
assign W_I_STAGE_LUT[281] = -16'd194;
assign W_R_STAGE_LUT[282] = 16'd166;
assign W_I_STAGE_LUT[282] = -16'd195;
assign W_R_STAGE_LUT[283] = 16'd165;
assign W_I_STAGE_LUT[283] = -16'd195;
assign W_R_STAGE_LUT[284] = 16'd165;
assign W_I_STAGE_LUT[284] = -16'd196;
assign W_R_STAGE_LUT[285] = 16'd164;
assign W_I_STAGE_LUT[285] = -16'd196;
assign W_R_STAGE_LUT[286] = 16'd164;
assign W_I_STAGE_LUT[286] = -16'd197;
assign W_R_STAGE_LUT[287] = 16'd163;
assign W_I_STAGE_LUT[287] = -16'd197;
assign W_R_STAGE_LUT[288] = 16'd162;
assign W_I_STAGE_LUT[288] = -16'd198;
assign W_R_STAGE_LUT[289] = 16'd162;
assign W_I_STAGE_LUT[289] = -16'd198;
assign W_R_STAGE_LUT[290] = 16'd161;
assign W_I_STAGE_LUT[290] = -16'd199;
assign W_R_STAGE_LUT[291] = 16'd161;
assign W_I_STAGE_LUT[291] = -16'd199;
assign W_R_STAGE_LUT[292] = 16'd160;
assign W_I_STAGE_LUT[292] = -16'd200;
assign W_R_STAGE_LUT[293] = 16'd159;
assign W_I_STAGE_LUT[293] = -16'd200;
assign W_R_STAGE_LUT[294] = 16'd159;
assign W_I_STAGE_LUT[294] = -16'd201;
assign W_R_STAGE_LUT[295] = 16'd158;
assign W_I_STAGE_LUT[295] = -16'd201;
assign W_R_STAGE_LUT[296] = 16'd157;
assign W_I_STAGE_LUT[296] = -16'd202;
assign W_R_STAGE_LUT[297] = 16'd157;
assign W_I_STAGE_LUT[297] = -16'd202;
assign W_R_STAGE_LUT[298] = 16'd156;
assign W_I_STAGE_LUT[298] = -16'd203;
assign W_R_STAGE_LUT[299] = 16'd156;
assign W_I_STAGE_LUT[299] = -16'd203;
assign W_R_STAGE_LUT[300] = 16'd155;
assign W_I_STAGE_LUT[300] = -16'd204;
assign W_R_STAGE_LUT[301] = 16'd154;
assign W_I_STAGE_LUT[301] = -16'd204;
assign W_R_STAGE_LUT[302] = 16'd154;
assign W_I_STAGE_LUT[302] = -16'd205;
assign W_R_STAGE_LUT[303] = 16'd153;
assign W_I_STAGE_LUT[303] = -16'd205;
assign W_R_STAGE_LUT[304] = 16'd152;
assign W_I_STAGE_LUT[304] = -16'd206;
assign W_R_STAGE_LUT[305] = 16'd152;
assign W_I_STAGE_LUT[305] = -16'd206;
assign W_R_STAGE_LUT[306] = 16'd151;
assign W_I_STAGE_LUT[306] = -16'd207;
assign W_R_STAGE_LUT[307] = 16'd151;
assign W_I_STAGE_LUT[307] = -16'd207;
assign W_R_STAGE_LUT[308] = 16'd150;
assign W_I_STAGE_LUT[308] = -16'd207;
assign W_R_STAGE_LUT[309] = 16'd149;
assign W_I_STAGE_LUT[309] = -16'd208;
assign W_R_STAGE_LUT[310] = 16'd149;
assign W_I_STAGE_LUT[310] = -16'd208;
assign W_R_STAGE_LUT[311] = 16'd148;
assign W_I_STAGE_LUT[311] = -16'd209;
assign W_R_STAGE_LUT[312] = 16'd147;
assign W_I_STAGE_LUT[312] = -16'd209;
assign W_R_STAGE_LUT[313] = 16'd147;
assign W_I_STAGE_LUT[313] = -16'd210;
assign W_R_STAGE_LUT[314] = 16'd146;
assign W_I_STAGE_LUT[314] = -16'd210;
assign W_R_STAGE_LUT[315] = 16'd145;
assign W_I_STAGE_LUT[315] = -16'd211;
assign W_R_STAGE_LUT[316] = 16'd145;
assign W_I_STAGE_LUT[316] = -16'd211;
assign W_R_STAGE_LUT[317] = 16'd144;
assign W_I_STAGE_LUT[317] = -16'd212;
assign W_R_STAGE_LUT[318] = 16'd144;
assign W_I_STAGE_LUT[318] = -16'd212;
assign W_R_STAGE_LUT[319] = 16'd143;
assign W_I_STAGE_LUT[319] = -16'd212;
assign W_R_STAGE_LUT[320] = 16'd142;
assign W_I_STAGE_LUT[320] = -16'd213;
assign W_R_STAGE_LUT[321] = 16'd142;
assign W_I_STAGE_LUT[321] = -16'd213;
assign W_R_STAGE_LUT[322] = 16'd141;
assign W_I_STAGE_LUT[322] = -16'd214;
assign W_R_STAGE_LUT[323] = 16'd140;
assign W_I_STAGE_LUT[323] = -16'd214;
assign W_R_STAGE_LUT[324] = 16'd140;
assign W_I_STAGE_LUT[324] = -16'd215;
assign W_R_STAGE_LUT[325] = 16'd139;
assign W_I_STAGE_LUT[325] = -16'd215;
assign W_R_STAGE_LUT[326] = 16'd138;
assign W_I_STAGE_LUT[326] = -16'd215;
assign W_R_STAGE_LUT[327] = 16'd138;
assign W_I_STAGE_LUT[327] = -16'd216;
assign W_R_STAGE_LUT[328] = 16'd137;
assign W_I_STAGE_LUT[328] = -16'd216;
assign W_R_STAGE_LUT[329] = 16'd136;
assign W_I_STAGE_LUT[329] = -16'd217;
assign W_R_STAGE_LUT[330] = 16'd136;
assign W_I_STAGE_LUT[330] = -16'd217;
assign W_R_STAGE_LUT[331] = 16'd135;
assign W_I_STAGE_LUT[331] = -16'd218;
assign W_R_STAGE_LUT[332] = 16'd134;
assign W_I_STAGE_LUT[332] = -16'd218;
assign W_R_STAGE_LUT[333] = 16'd134;
assign W_I_STAGE_LUT[333] = -16'd218;
assign W_R_STAGE_LUT[334] = 16'd133;
assign W_I_STAGE_LUT[334] = -16'd219;
assign W_R_STAGE_LUT[335] = 16'd132;
assign W_I_STAGE_LUT[335] = -16'd219;
assign W_R_STAGE_LUT[336] = 16'd132;
assign W_I_STAGE_LUT[336] = -16'd220;
assign W_R_STAGE_LUT[337] = 16'd131;
assign W_I_STAGE_LUT[337] = -16'd220;
assign W_R_STAGE_LUT[338] = 16'd130;
assign W_I_STAGE_LUT[338] = -16'd220;
assign W_R_STAGE_LUT[339] = 16'd130;
assign W_I_STAGE_LUT[339] = -16'd221;
assign W_R_STAGE_LUT[340] = 16'd129;
assign W_I_STAGE_LUT[340] = -16'd221;
assign W_R_STAGE_LUT[341] = 16'd128;
assign W_I_STAGE_LUT[341] = -16'd222;
assign W_R_STAGE_LUT[342] = 16'd128;
assign W_I_STAGE_LUT[342] = -16'd222;
assign W_R_STAGE_LUT[343] = 16'd127;
assign W_I_STAGE_LUT[343] = -16'd222;
assign W_R_STAGE_LUT[344] = 16'd126;
assign W_I_STAGE_LUT[344] = -16'd223;
assign W_R_STAGE_LUT[345] = 16'd125;
assign W_I_STAGE_LUT[345] = -16'd223;
assign W_R_STAGE_LUT[346] = 16'd125;
assign W_I_STAGE_LUT[346] = -16'd224;
assign W_R_STAGE_LUT[347] = 16'd124;
assign W_I_STAGE_LUT[347] = -16'd224;
assign W_R_STAGE_LUT[348] = 16'd123;
assign W_I_STAGE_LUT[348] = -16'd224;
assign W_R_STAGE_LUT[349] = 16'd123;
assign W_I_STAGE_LUT[349] = -16'd225;
assign W_R_STAGE_LUT[350] = 16'd122;
assign W_I_STAGE_LUT[350] = -16'd225;
assign W_R_STAGE_LUT[351] = 16'd121;
assign W_I_STAGE_LUT[351] = -16'd225;
assign W_R_STAGE_LUT[352] = 16'd121;
assign W_I_STAGE_LUT[352] = -16'd226;
assign W_R_STAGE_LUT[353] = 16'd120;
assign W_I_STAGE_LUT[353] = -16'd226;
assign W_R_STAGE_LUT[354] = 16'd119;
assign W_I_STAGE_LUT[354] = -16'd227;
assign W_R_STAGE_LUT[355] = 16'd119;
assign W_I_STAGE_LUT[355] = -16'd227;
assign W_R_STAGE_LUT[356] = 16'd118;
assign W_I_STAGE_LUT[356] = -16'd227;
assign W_R_STAGE_LUT[357] = 16'd117;
assign W_I_STAGE_LUT[357] = -16'd228;
assign W_R_STAGE_LUT[358] = 16'd117;
assign W_I_STAGE_LUT[358] = -16'd228;
assign W_R_STAGE_LUT[359] = 16'd116;
assign W_I_STAGE_LUT[359] = -16'd228;
assign W_R_STAGE_LUT[360] = 16'd115;
assign W_I_STAGE_LUT[360] = -16'd229;
assign W_R_STAGE_LUT[361] = 16'd114;
assign W_I_STAGE_LUT[361] = -16'd229;
assign W_R_STAGE_LUT[362] = 16'd114;
assign W_I_STAGE_LUT[362] = -16'd229;
assign W_R_STAGE_LUT[363] = 16'd113;
assign W_I_STAGE_LUT[363] = -16'd230;
assign W_R_STAGE_LUT[364] = 16'd112;
assign W_I_STAGE_LUT[364] = -16'd230;
assign W_R_STAGE_LUT[365] = 16'd112;
assign W_I_STAGE_LUT[365] = -16'd230;
assign W_R_STAGE_LUT[366] = 16'd111;
assign W_I_STAGE_LUT[366] = -16'd231;
assign W_R_STAGE_LUT[367] = 16'd110;
assign W_I_STAGE_LUT[367] = -16'd231;
assign W_R_STAGE_LUT[368] = 16'd109;
assign W_I_STAGE_LUT[368] = -16'd231;
assign W_R_STAGE_LUT[369] = 16'd109;
assign W_I_STAGE_LUT[369] = -16'd232;
assign W_R_STAGE_LUT[370] = 16'd108;
assign W_I_STAGE_LUT[370] = -16'd232;
assign W_R_STAGE_LUT[371] = 16'd107;
assign W_I_STAGE_LUT[371] = -16'd232;
assign W_R_STAGE_LUT[372] = 16'd107;
assign W_I_STAGE_LUT[372] = -16'd233;
assign W_R_STAGE_LUT[373] = 16'd106;
assign W_I_STAGE_LUT[373] = -16'd233;
assign W_R_STAGE_LUT[374] = 16'd105;
assign W_I_STAGE_LUT[374] = -16'd233;
assign W_R_STAGE_LUT[375] = 16'd104;
assign W_I_STAGE_LUT[375] = -16'd234;
assign W_R_STAGE_LUT[376] = 16'd104;
assign W_I_STAGE_LUT[376] = -16'd234;
assign W_R_STAGE_LUT[377] = 16'd103;
assign W_I_STAGE_LUT[377] = -16'd234;
assign W_R_STAGE_LUT[378] = 16'd102;
assign W_I_STAGE_LUT[378] = -16'd235;
assign W_R_STAGE_LUT[379] = 16'd102;
assign W_I_STAGE_LUT[379] = -16'd235;
assign W_R_STAGE_LUT[380] = 16'd101;
assign W_I_STAGE_LUT[380] = -16'd235;
assign W_R_STAGE_LUT[381] = 16'd100;
assign W_I_STAGE_LUT[381] = -16'd236;
assign W_R_STAGE_LUT[382] = 16'd99;
assign W_I_STAGE_LUT[382] = -16'd236;
assign W_R_STAGE_LUT[383] = 16'd99;
assign W_I_STAGE_LUT[383] = -16'd236;
assign W_R_STAGE_LUT[384] = 16'd98;
assign W_I_STAGE_LUT[384] = -16'd237;
assign W_R_STAGE_LUT[385] = 16'd97;
assign W_I_STAGE_LUT[385] = -16'd237;
assign W_R_STAGE_LUT[386] = 16'd97;
assign W_I_STAGE_LUT[386] = -16'd237;
assign W_R_STAGE_LUT[387] = 16'd96;
assign W_I_STAGE_LUT[387] = -16'd237;
assign W_R_STAGE_LUT[388] = 16'd95;
assign W_I_STAGE_LUT[388] = -16'd238;
assign W_R_STAGE_LUT[389] = 16'd94;
assign W_I_STAGE_LUT[389] = -16'd238;
assign W_R_STAGE_LUT[390] = 16'd94;
assign W_I_STAGE_LUT[390] = -16'd238;
assign W_R_STAGE_LUT[391] = 16'd93;
assign W_I_STAGE_LUT[391] = -16'd239;
assign W_R_STAGE_LUT[392] = 16'd92;
assign W_I_STAGE_LUT[392] = -16'd239;
assign W_R_STAGE_LUT[393] = 16'd91;
assign W_I_STAGE_LUT[393] = -16'd239;
assign W_R_STAGE_LUT[394] = 16'd91;
assign W_I_STAGE_LUT[394] = -16'd239;
assign W_R_STAGE_LUT[395] = 16'd90;
assign W_I_STAGE_LUT[395] = -16'd240;
assign W_R_STAGE_LUT[396] = 16'd89;
assign W_I_STAGE_LUT[396] = -16'd240;
assign W_R_STAGE_LUT[397] = 16'd88;
assign W_I_STAGE_LUT[397] = -16'd240;
assign W_R_STAGE_LUT[398] = 16'd88;
assign W_I_STAGE_LUT[398] = -16'd241;
assign W_R_STAGE_LUT[399] = 16'd87;
assign W_I_STAGE_LUT[399] = -16'd241;
assign W_R_STAGE_LUT[400] = 16'd86;
assign W_I_STAGE_LUT[400] = -16'd241;
assign W_R_STAGE_LUT[401] = 16'd86;
assign W_I_STAGE_LUT[401] = -16'd241;
assign W_R_STAGE_LUT[402] = 16'd85;
assign W_I_STAGE_LUT[402] = -16'd242;
assign W_R_STAGE_LUT[403] = 16'd84;
assign W_I_STAGE_LUT[403] = -16'd242;
assign W_R_STAGE_LUT[404] = 16'd83;
assign W_I_STAGE_LUT[404] = -16'd242;
assign W_R_STAGE_LUT[405] = 16'd83;
assign W_I_STAGE_LUT[405] = -16'd242;
assign W_R_STAGE_LUT[406] = 16'd82;
assign W_I_STAGE_LUT[406] = -16'd243;
assign W_R_STAGE_LUT[407] = 16'd81;
assign W_I_STAGE_LUT[407] = -16'd243;
assign W_R_STAGE_LUT[408] = 16'd80;
assign W_I_STAGE_LUT[408] = -16'd243;
assign W_R_STAGE_LUT[409] = 16'd80;
assign W_I_STAGE_LUT[409] = -16'd243;
assign W_R_STAGE_LUT[410] = 16'd79;
assign W_I_STAGE_LUT[410] = -16'd244;
assign W_R_STAGE_LUT[411] = 16'd78;
assign W_I_STAGE_LUT[411] = -16'd244;
assign W_R_STAGE_LUT[412] = 16'd77;
assign W_I_STAGE_LUT[412] = -16'd244;
assign W_R_STAGE_LUT[413] = 16'd77;
assign W_I_STAGE_LUT[413] = -16'd244;
assign W_R_STAGE_LUT[414] = 16'd76;
assign W_I_STAGE_LUT[414] = -16'd245;
assign W_R_STAGE_LUT[415] = 16'd75;
assign W_I_STAGE_LUT[415] = -16'd245;
assign W_R_STAGE_LUT[416] = 16'd74;
assign W_I_STAGE_LUT[416] = -16'd245;
assign W_R_STAGE_LUT[417] = 16'd74;
assign W_I_STAGE_LUT[417] = -16'd245;
assign W_R_STAGE_LUT[418] = 16'd73;
assign W_I_STAGE_LUT[418] = -16'd245;
assign W_R_STAGE_LUT[419] = 16'd72;
assign W_I_STAGE_LUT[419] = -16'd246;
assign W_R_STAGE_LUT[420] = 16'd71;
assign W_I_STAGE_LUT[420] = -16'd246;
assign W_R_STAGE_LUT[421] = 16'd71;
assign W_I_STAGE_LUT[421] = -16'd246;
assign W_R_STAGE_LUT[422] = 16'd70;
assign W_I_STAGE_LUT[422] = -16'd246;
assign W_R_STAGE_LUT[423] = 16'd69;
assign W_I_STAGE_LUT[423] = -16'd247;
assign W_R_STAGE_LUT[424] = 16'd68;
assign W_I_STAGE_LUT[424] = -16'd247;
assign W_R_STAGE_LUT[425] = 16'd68;
assign W_I_STAGE_LUT[425] = -16'd247;
assign W_R_STAGE_LUT[426] = 16'd67;
assign W_I_STAGE_LUT[426] = -16'd247;
assign W_R_STAGE_LUT[427] = 16'd66;
assign W_I_STAGE_LUT[427] = -16'd247;
assign W_R_STAGE_LUT[428] = 16'd65;
assign W_I_STAGE_LUT[428] = -16'd248;
assign W_R_STAGE_LUT[429] = 16'd64;
assign W_I_STAGE_LUT[429] = -16'd248;
assign W_R_STAGE_LUT[430] = 16'd64;
assign W_I_STAGE_LUT[430] = -16'd248;
assign W_R_STAGE_LUT[431] = 16'd63;
assign W_I_STAGE_LUT[431] = -16'd248;
assign W_R_STAGE_LUT[432] = 16'd62;
assign W_I_STAGE_LUT[432] = -16'd248;
assign W_R_STAGE_LUT[433] = 16'd61;
assign W_I_STAGE_LUT[433] = -16'd249;
assign W_R_STAGE_LUT[434] = 16'd61;
assign W_I_STAGE_LUT[434] = -16'd249;
assign W_R_STAGE_LUT[435] = 16'd60;
assign W_I_STAGE_LUT[435] = -16'd249;
assign W_R_STAGE_LUT[436] = 16'd59;
assign W_I_STAGE_LUT[436] = -16'd249;
assign W_R_STAGE_LUT[437] = 16'd58;
assign W_I_STAGE_LUT[437] = -16'd249;
assign W_R_STAGE_LUT[438] = 16'd58;
assign W_I_STAGE_LUT[438] = -16'd249;
assign W_R_STAGE_LUT[439] = 16'd57;
assign W_I_STAGE_LUT[439] = -16'd250;
assign W_R_STAGE_LUT[440] = 16'd56;
assign W_I_STAGE_LUT[440] = -16'd250;
assign W_R_STAGE_LUT[441] = 16'd55;
assign W_I_STAGE_LUT[441] = -16'd250;
assign W_R_STAGE_LUT[442] = 16'd55;
assign W_I_STAGE_LUT[442] = -16'd250;
assign W_R_STAGE_LUT[443] = 16'd54;
assign W_I_STAGE_LUT[443] = -16'd250;
assign W_R_STAGE_LUT[444] = 16'd53;
assign W_I_STAGE_LUT[444] = -16'd250;
assign W_R_STAGE_LUT[445] = 16'd52;
assign W_I_STAGE_LUT[445] = -16'd251;
assign W_R_STAGE_LUT[446] = 16'd51;
assign W_I_STAGE_LUT[446] = -16'd251;
assign W_R_STAGE_LUT[447] = 16'd51;
assign W_I_STAGE_LUT[447] = -16'd251;
assign W_R_STAGE_LUT[448] = 16'd50;
assign W_I_STAGE_LUT[448] = -16'd251;
assign W_R_STAGE_LUT[449] = 16'd49;
assign W_I_STAGE_LUT[449] = -16'd251;
assign W_R_STAGE_LUT[450] = 16'd48;
assign W_I_STAGE_LUT[450] = -16'd251;
assign W_R_STAGE_LUT[451] = 16'd48;
assign W_I_STAGE_LUT[451] = -16'd252;
assign W_R_STAGE_LUT[452] = 16'd47;
assign W_I_STAGE_LUT[452] = -16'd252;
assign W_R_STAGE_LUT[453] = 16'd46;
assign W_I_STAGE_LUT[453] = -16'd252;
assign W_R_STAGE_LUT[454] = 16'd45;
assign W_I_STAGE_LUT[454] = -16'd252;
assign W_R_STAGE_LUT[455] = 16'd45;
assign W_I_STAGE_LUT[455] = -16'd252;
assign W_R_STAGE_LUT[456] = 16'd44;
assign W_I_STAGE_LUT[456] = -16'd252;
assign W_R_STAGE_LUT[457] = 16'd43;
assign W_I_STAGE_LUT[457] = -16'd252;
assign W_R_STAGE_LUT[458] = 16'd42;
assign W_I_STAGE_LUT[458] = -16'd252;
assign W_R_STAGE_LUT[459] = 16'd41;
assign W_I_STAGE_LUT[459] = -16'd253;
assign W_R_STAGE_LUT[460] = 16'd41;
assign W_I_STAGE_LUT[460] = -16'd253;
assign W_R_STAGE_LUT[461] = 16'd40;
assign W_I_STAGE_LUT[461] = -16'd253;
assign W_R_STAGE_LUT[462] = 16'd39;
assign W_I_STAGE_LUT[462] = -16'd253;
assign W_R_STAGE_LUT[463] = 16'd38;
assign W_I_STAGE_LUT[463] = -16'd253;
assign W_R_STAGE_LUT[464] = 16'd38;
assign W_I_STAGE_LUT[464] = -16'd253;
assign W_R_STAGE_LUT[465] = 16'd37;
assign W_I_STAGE_LUT[465] = -16'd253;
assign W_R_STAGE_LUT[466] = 16'd36;
assign W_I_STAGE_LUT[466] = -16'd253;
assign W_R_STAGE_LUT[467] = 16'd35;
assign W_I_STAGE_LUT[467] = -16'd254;
assign W_R_STAGE_LUT[468] = 16'd34;
assign W_I_STAGE_LUT[468] = -16'd254;
assign W_R_STAGE_LUT[469] = 16'd34;
assign W_I_STAGE_LUT[469] = -16'd254;
assign W_R_STAGE_LUT[470] = 16'd33;
assign W_I_STAGE_LUT[470] = -16'd254;
assign W_R_STAGE_LUT[471] = 16'd32;
assign W_I_STAGE_LUT[471] = -16'd254;
assign W_R_STAGE_LUT[472] = 16'd31;
assign W_I_STAGE_LUT[472] = -16'd254;
assign W_R_STAGE_LUT[473] = 16'd31;
assign W_I_STAGE_LUT[473] = -16'd254;
assign W_R_STAGE_LUT[474] = 16'd30;
assign W_I_STAGE_LUT[474] = -16'd254;
assign W_R_STAGE_LUT[475] = 16'd29;
assign W_I_STAGE_LUT[475] = -16'd254;
assign W_R_STAGE_LUT[476] = 16'd28;
assign W_I_STAGE_LUT[476] = -16'd254;
assign W_R_STAGE_LUT[477] = 16'd27;
assign W_I_STAGE_LUT[477] = -16'd255;
assign W_R_STAGE_LUT[478] = 16'd27;
assign W_I_STAGE_LUT[478] = -16'd255;
assign W_R_STAGE_LUT[479] = 16'd26;
assign W_I_STAGE_LUT[479] = -16'd255;
assign W_R_STAGE_LUT[480] = 16'd25;
assign W_I_STAGE_LUT[480] = -16'd255;
assign W_R_STAGE_LUT[481] = 16'd24;
assign W_I_STAGE_LUT[481] = -16'd255;
assign W_R_STAGE_LUT[482] = 16'd24;
assign W_I_STAGE_LUT[482] = -16'd255;
assign W_R_STAGE_LUT[483] = 16'd23;
assign W_I_STAGE_LUT[483] = -16'd255;
assign W_R_STAGE_LUT[484] = 16'd22;
assign W_I_STAGE_LUT[484] = -16'd255;
assign W_R_STAGE_LUT[485] = 16'd21;
assign W_I_STAGE_LUT[485] = -16'd255;
assign W_R_STAGE_LUT[486] = 16'd20;
assign W_I_STAGE_LUT[486] = -16'd255;
assign W_R_STAGE_LUT[487] = 16'd20;
assign W_I_STAGE_LUT[487] = -16'd255;
assign W_R_STAGE_LUT[488] = 16'd19;
assign W_I_STAGE_LUT[488] = -16'd255;
assign W_R_STAGE_LUT[489] = 16'd18;
assign W_I_STAGE_LUT[489] = -16'd255;
assign W_R_STAGE_LUT[490] = 16'd17;
assign W_I_STAGE_LUT[490] = -16'd255;
assign W_R_STAGE_LUT[491] = 16'd16;
assign W_I_STAGE_LUT[491] = -16'd255;
assign W_R_STAGE_LUT[492] = 16'd16;
assign W_I_STAGE_LUT[492] = -16'd256;
assign W_R_STAGE_LUT[493] = 16'd15;
assign W_I_STAGE_LUT[493] = -16'd256;
assign W_R_STAGE_LUT[494] = 16'd14;
assign W_I_STAGE_LUT[494] = -16'd256;
assign W_R_STAGE_LUT[495] = 16'd13;
assign W_I_STAGE_LUT[495] = -16'd256;
assign W_R_STAGE_LUT[496] = 16'd13;
assign W_I_STAGE_LUT[496] = -16'd256;
assign W_R_STAGE_LUT[497] = 16'd12;
assign W_I_STAGE_LUT[497] = -16'd256;
assign W_R_STAGE_LUT[498] = 16'd11;
assign W_I_STAGE_LUT[498] = -16'd256;
assign W_R_STAGE_LUT[499] = 16'd10;
assign W_I_STAGE_LUT[499] = -16'd256;
assign W_R_STAGE_LUT[500] = 16'd9;
assign W_I_STAGE_LUT[500] = -16'd256;
assign W_R_STAGE_LUT[501] = 16'd9;
assign W_I_STAGE_LUT[501] = -16'd256;
assign W_R_STAGE_LUT[502] = 16'd8;
assign W_I_STAGE_LUT[502] = -16'd256;
assign W_R_STAGE_LUT[503] = 16'd7;
assign W_I_STAGE_LUT[503] = -16'd256;
assign W_R_STAGE_LUT[504] = 16'd6;
assign W_I_STAGE_LUT[504] = -16'd256;
assign W_R_STAGE_LUT[505] = 16'd5;
assign W_I_STAGE_LUT[505] = -16'd256;
assign W_R_STAGE_LUT[506] = 16'd5;
assign W_I_STAGE_LUT[506] = -16'd256;
assign W_R_STAGE_LUT[507] = 16'd4;
assign W_I_STAGE_LUT[507] = -16'd256;
assign W_R_STAGE_LUT[508] = 16'd3;
assign W_I_STAGE_LUT[508] = -16'd256;
assign W_R_STAGE_LUT[509] = 16'd2;
assign W_I_STAGE_LUT[509] = -16'd256;
assign W_R_STAGE_LUT[510] = 16'd2;
assign W_I_STAGE_LUT[510] = -16'd256;
assign W_R_STAGE_LUT[511] = 16'd1;
assign W_I_STAGE_LUT[511] = -16'd256;
assign W_R_STAGE_LUT[512] = 16'd0;
assign W_I_STAGE_LUT[512] = -16'd256;
assign W_R_STAGE_LUT[513] = -16'd1;
assign W_I_STAGE_LUT[513] = -16'd256;
assign W_R_STAGE_LUT[514] = -16'd2;
assign W_I_STAGE_LUT[514] = -16'd256;
assign W_R_STAGE_LUT[515] = -16'd2;
assign W_I_STAGE_LUT[515] = -16'd256;
assign W_R_STAGE_LUT[516] = -16'd3;
assign W_I_STAGE_LUT[516] = -16'd256;
assign W_R_STAGE_LUT[517] = -16'd4;
assign W_I_STAGE_LUT[517] = -16'd256;
assign W_R_STAGE_LUT[518] = -16'd5;
assign W_I_STAGE_LUT[518] = -16'd256;
assign W_R_STAGE_LUT[519] = -16'd5;
assign W_I_STAGE_LUT[519] = -16'd256;
assign W_R_STAGE_LUT[520] = -16'd6;
assign W_I_STAGE_LUT[520] = -16'd256;
assign W_R_STAGE_LUT[521] = -16'd7;
assign W_I_STAGE_LUT[521] = -16'd256;
assign W_R_STAGE_LUT[522] = -16'd8;
assign W_I_STAGE_LUT[522] = -16'd256;
assign W_R_STAGE_LUT[523] = -16'd9;
assign W_I_STAGE_LUT[523] = -16'd256;
assign W_R_STAGE_LUT[524] = -16'd9;
assign W_I_STAGE_LUT[524] = -16'd256;
assign W_R_STAGE_LUT[525] = -16'd10;
assign W_I_STAGE_LUT[525] = -16'd256;
assign W_R_STAGE_LUT[526] = -16'd11;
assign W_I_STAGE_LUT[526] = -16'd256;
assign W_R_STAGE_LUT[527] = -16'd12;
assign W_I_STAGE_LUT[527] = -16'd256;
assign W_R_STAGE_LUT[528] = -16'd13;
assign W_I_STAGE_LUT[528] = -16'd256;
assign W_R_STAGE_LUT[529] = -16'd13;
assign W_I_STAGE_LUT[529] = -16'd256;
assign W_R_STAGE_LUT[530] = -16'd14;
assign W_I_STAGE_LUT[530] = -16'd256;
assign W_R_STAGE_LUT[531] = -16'd15;
assign W_I_STAGE_LUT[531] = -16'd256;
assign W_R_STAGE_LUT[532] = -16'd16;
assign W_I_STAGE_LUT[532] = -16'd256;
assign W_R_STAGE_LUT[533] = -16'd16;
assign W_I_STAGE_LUT[533] = -16'd255;
assign W_R_STAGE_LUT[534] = -16'd17;
assign W_I_STAGE_LUT[534] = -16'd255;
assign W_R_STAGE_LUT[535] = -16'd18;
assign W_I_STAGE_LUT[535] = -16'd255;
assign W_R_STAGE_LUT[536] = -16'd19;
assign W_I_STAGE_LUT[536] = -16'd255;
assign W_R_STAGE_LUT[537] = -16'd20;
assign W_I_STAGE_LUT[537] = -16'd255;
assign W_R_STAGE_LUT[538] = -16'd20;
assign W_I_STAGE_LUT[538] = -16'd255;
assign W_R_STAGE_LUT[539] = -16'd21;
assign W_I_STAGE_LUT[539] = -16'd255;
assign W_R_STAGE_LUT[540] = -16'd22;
assign W_I_STAGE_LUT[540] = -16'd255;
assign W_R_STAGE_LUT[541] = -16'd23;
assign W_I_STAGE_LUT[541] = -16'd255;
assign W_R_STAGE_LUT[542] = -16'd24;
assign W_I_STAGE_LUT[542] = -16'd255;
assign W_R_STAGE_LUT[543] = -16'd24;
assign W_I_STAGE_LUT[543] = -16'd255;
assign W_R_STAGE_LUT[544] = -16'd25;
assign W_I_STAGE_LUT[544] = -16'd255;
assign W_R_STAGE_LUT[545] = -16'd26;
assign W_I_STAGE_LUT[545] = -16'd255;
assign W_R_STAGE_LUT[546] = -16'd27;
assign W_I_STAGE_LUT[546] = -16'd255;
assign W_R_STAGE_LUT[547] = -16'd27;
assign W_I_STAGE_LUT[547] = -16'd255;
assign W_R_STAGE_LUT[548] = -16'd28;
assign W_I_STAGE_LUT[548] = -16'd254;
assign W_R_STAGE_LUT[549] = -16'd29;
assign W_I_STAGE_LUT[549] = -16'd254;
assign W_R_STAGE_LUT[550] = -16'd30;
assign W_I_STAGE_LUT[550] = -16'd254;
assign W_R_STAGE_LUT[551] = -16'd31;
assign W_I_STAGE_LUT[551] = -16'd254;
assign W_R_STAGE_LUT[552] = -16'd31;
assign W_I_STAGE_LUT[552] = -16'd254;
assign W_R_STAGE_LUT[553] = -16'd32;
assign W_I_STAGE_LUT[553] = -16'd254;
assign W_R_STAGE_LUT[554] = -16'd33;
assign W_I_STAGE_LUT[554] = -16'd254;
assign W_R_STAGE_LUT[555] = -16'd34;
assign W_I_STAGE_LUT[555] = -16'd254;
assign W_R_STAGE_LUT[556] = -16'd34;
assign W_I_STAGE_LUT[556] = -16'd254;
assign W_R_STAGE_LUT[557] = -16'd35;
assign W_I_STAGE_LUT[557] = -16'd254;
assign W_R_STAGE_LUT[558] = -16'd36;
assign W_I_STAGE_LUT[558] = -16'd253;
assign W_R_STAGE_LUT[559] = -16'd37;
assign W_I_STAGE_LUT[559] = -16'd253;
assign W_R_STAGE_LUT[560] = -16'd38;
assign W_I_STAGE_LUT[560] = -16'd253;
assign W_R_STAGE_LUT[561] = -16'd38;
assign W_I_STAGE_LUT[561] = -16'd253;
assign W_R_STAGE_LUT[562] = -16'd39;
assign W_I_STAGE_LUT[562] = -16'd253;
assign W_R_STAGE_LUT[563] = -16'd40;
assign W_I_STAGE_LUT[563] = -16'd253;
assign W_R_STAGE_LUT[564] = -16'd41;
assign W_I_STAGE_LUT[564] = -16'd253;
assign W_R_STAGE_LUT[565] = -16'd41;
assign W_I_STAGE_LUT[565] = -16'd253;
assign W_R_STAGE_LUT[566] = -16'd42;
assign W_I_STAGE_LUT[566] = -16'd252;
assign W_R_STAGE_LUT[567] = -16'd43;
assign W_I_STAGE_LUT[567] = -16'd252;
assign W_R_STAGE_LUT[568] = -16'd44;
assign W_I_STAGE_LUT[568] = -16'd252;
assign W_R_STAGE_LUT[569] = -16'd45;
assign W_I_STAGE_LUT[569] = -16'd252;
assign W_R_STAGE_LUT[570] = -16'd45;
assign W_I_STAGE_LUT[570] = -16'd252;
assign W_R_STAGE_LUT[571] = -16'd46;
assign W_I_STAGE_LUT[571] = -16'd252;
assign W_R_STAGE_LUT[572] = -16'd47;
assign W_I_STAGE_LUT[572] = -16'd252;
assign W_R_STAGE_LUT[573] = -16'd48;
assign W_I_STAGE_LUT[573] = -16'd252;
assign W_R_STAGE_LUT[574] = -16'd48;
assign W_I_STAGE_LUT[574] = -16'd251;
assign W_R_STAGE_LUT[575] = -16'd49;
assign W_I_STAGE_LUT[575] = -16'd251;
assign W_R_STAGE_LUT[576] = -16'd50;
assign W_I_STAGE_LUT[576] = -16'd251;
assign W_R_STAGE_LUT[577] = -16'd51;
assign W_I_STAGE_LUT[577] = -16'd251;
assign W_R_STAGE_LUT[578] = -16'd51;
assign W_I_STAGE_LUT[578] = -16'd251;
assign W_R_STAGE_LUT[579] = -16'd52;
assign W_I_STAGE_LUT[579] = -16'd251;
assign W_R_STAGE_LUT[580] = -16'd53;
assign W_I_STAGE_LUT[580] = -16'd250;
assign W_R_STAGE_LUT[581] = -16'd54;
assign W_I_STAGE_LUT[581] = -16'd250;
assign W_R_STAGE_LUT[582] = -16'd55;
assign W_I_STAGE_LUT[582] = -16'd250;
assign W_R_STAGE_LUT[583] = -16'd55;
assign W_I_STAGE_LUT[583] = -16'd250;
assign W_R_STAGE_LUT[584] = -16'd56;
assign W_I_STAGE_LUT[584] = -16'd250;
assign W_R_STAGE_LUT[585] = -16'd57;
assign W_I_STAGE_LUT[585] = -16'd250;
assign W_R_STAGE_LUT[586] = -16'd58;
assign W_I_STAGE_LUT[586] = -16'd249;
assign W_R_STAGE_LUT[587] = -16'd58;
assign W_I_STAGE_LUT[587] = -16'd249;
assign W_R_STAGE_LUT[588] = -16'd59;
assign W_I_STAGE_LUT[588] = -16'd249;
assign W_R_STAGE_LUT[589] = -16'd60;
assign W_I_STAGE_LUT[589] = -16'd249;
assign W_R_STAGE_LUT[590] = -16'd61;
assign W_I_STAGE_LUT[590] = -16'd249;
assign W_R_STAGE_LUT[591] = -16'd61;
assign W_I_STAGE_LUT[591] = -16'd249;
assign W_R_STAGE_LUT[592] = -16'd62;
assign W_I_STAGE_LUT[592] = -16'd248;
assign W_R_STAGE_LUT[593] = -16'd63;
assign W_I_STAGE_LUT[593] = -16'd248;
assign W_R_STAGE_LUT[594] = -16'd64;
assign W_I_STAGE_LUT[594] = -16'd248;
assign W_R_STAGE_LUT[595] = -16'd64;
assign W_I_STAGE_LUT[595] = -16'd248;
assign W_R_STAGE_LUT[596] = -16'd65;
assign W_I_STAGE_LUT[596] = -16'd248;
assign W_R_STAGE_LUT[597] = -16'd66;
assign W_I_STAGE_LUT[597] = -16'd247;
assign W_R_STAGE_LUT[598] = -16'd67;
assign W_I_STAGE_LUT[598] = -16'd247;
assign W_R_STAGE_LUT[599] = -16'd68;
assign W_I_STAGE_LUT[599] = -16'd247;
assign W_R_STAGE_LUT[600] = -16'd68;
assign W_I_STAGE_LUT[600] = -16'd247;
assign W_R_STAGE_LUT[601] = -16'd69;
assign W_I_STAGE_LUT[601] = -16'd247;
assign W_R_STAGE_LUT[602] = -16'd70;
assign W_I_STAGE_LUT[602] = -16'd246;
assign W_R_STAGE_LUT[603] = -16'd71;
assign W_I_STAGE_LUT[603] = -16'd246;
assign W_R_STAGE_LUT[604] = -16'd71;
assign W_I_STAGE_LUT[604] = -16'd246;
assign W_R_STAGE_LUT[605] = -16'd72;
assign W_I_STAGE_LUT[605] = -16'd246;
assign W_R_STAGE_LUT[606] = -16'd73;
assign W_I_STAGE_LUT[606] = -16'd245;
assign W_R_STAGE_LUT[607] = -16'd74;
assign W_I_STAGE_LUT[607] = -16'd245;
assign W_R_STAGE_LUT[608] = -16'd74;
assign W_I_STAGE_LUT[608] = -16'd245;
assign W_R_STAGE_LUT[609] = -16'd75;
assign W_I_STAGE_LUT[609] = -16'd245;
assign W_R_STAGE_LUT[610] = -16'd76;
assign W_I_STAGE_LUT[610] = -16'd245;
assign W_R_STAGE_LUT[611] = -16'd77;
assign W_I_STAGE_LUT[611] = -16'd244;
assign W_R_STAGE_LUT[612] = -16'd77;
assign W_I_STAGE_LUT[612] = -16'd244;
assign W_R_STAGE_LUT[613] = -16'd78;
assign W_I_STAGE_LUT[613] = -16'd244;
assign W_R_STAGE_LUT[614] = -16'd79;
assign W_I_STAGE_LUT[614] = -16'd244;
assign W_R_STAGE_LUT[615] = -16'd80;
assign W_I_STAGE_LUT[615] = -16'd243;
assign W_R_STAGE_LUT[616] = -16'd80;
assign W_I_STAGE_LUT[616] = -16'd243;
assign W_R_STAGE_LUT[617] = -16'd81;
assign W_I_STAGE_LUT[617] = -16'd243;
assign W_R_STAGE_LUT[618] = -16'd82;
assign W_I_STAGE_LUT[618] = -16'd243;
assign W_R_STAGE_LUT[619] = -16'd83;
assign W_I_STAGE_LUT[619] = -16'd242;
assign W_R_STAGE_LUT[620] = -16'd83;
assign W_I_STAGE_LUT[620] = -16'd242;
assign W_R_STAGE_LUT[621] = -16'd84;
assign W_I_STAGE_LUT[621] = -16'd242;
assign W_R_STAGE_LUT[622] = -16'd85;
assign W_I_STAGE_LUT[622] = -16'd242;
assign W_R_STAGE_LUT[623] = -16'd86;
assign W_I_STAGE_LUT[623] = -16'd241;
assign W_R_STAGE_LUT[624] = -16'd86;
assign W_I_STAGE_LUT[624] = -16'd241;
assign W_R_STAGE_LUT[625] = -16'd87;
assign W_I_STAGE_LUT[625] = -16'd241;
assign W_R_STAGE_LUT[626] = -16'd88;
assign W_I_STAGE_LUT[626] = -16'd241;
assign W_R_STAGE_LUT[627] = -16'd88;
assign W_I_STAGE_LUT[627] = -16'd240;
assign W_R_STAGE_LUT[628] = -16'd89;
assign W_I_STAGE_LUT[628] = -16'd240;
assign W_R_STAGE_LUT[629] = -16'd90;
assign W_I_STAGE_LUT[629] = -16'd240;
assign W_R_STAGE_LUT[630] = -16'd91;
assign W_I_STAGE_LUT[630] = -16'd239;
assign W_R_STAGE_LUT[631] = -16'd91;
assign W_I_STAGE_LUT[631] = -16'd239;
assign W_R_STAGE_LUT[632] = -16'd92;
assign W_I_STAGE_LUT[632] = -16'd239;
assign W_R_STAGE_LUT[633] = -16'd93;
assign W_I_STAGE_LUT[633] = -16'd239;
assign W_R_STAGE_LUT[634] = -16'd94;
assign W_I_STAGE_LUT[634] = -16'd238;
assign W_R_STAGE_LUT[635] = -16'd94;
assign W_I_STAGE_LUT[635] = -16'd238;
assign W_R_STAGE_LUT[636] = -16'd95;
assign W_I_STAGE_LUT[636] = -16'd238;
assign W_R_STAGE_LUT[637] = -16'd96;
assign W_I_STAGE_LUT[637] = -16'd237;
assign W_R_STAGE_LUT[638] = -16'd97;
assign W_I_STAGE_LUT[638] = -16'd237;
assign W_R_STAGE_LUT[639] = -16'd97;
assign W_I_STAGE_LUT[639] = -16'd237;
assign W_R_STAGE_LUT[640] = -16'd98;
assign W_I_STAGE_LUT[640] = -16'd237;
assign W_R_STAGE_LUT[641] = -16'd99;
assign W_I_STAGE_LUT[641] = -16'd236;
assign W_R_STAGE_LUT[642] = -16'd99;
assign W_I_STAGE_LUT[642] = -16'd236;
assign W_R_STAGE_LUT[643] = -16'd100;
assign W_I_STAGE_LUT[643] = -16'd236;
assign W_R_STAGE_LUT[644] = -16'd101;
assign W_I_STAGE_LUT[644] = -16'd235;
assign W_R_STAGE_LUT[645] = -16'd102;
assign W_I_STAGE_LUT[645] = -16'd235;
assign W_R_STAGE_LUT[646] = -16'd102;
assign W_I_STAGE_LUT[646] = -16'd235;
assign W_R_STAGE_LUT[647] = -16'd103;
assign W_I_STAGE_LUT[647] = -16'd234;
assign W_R_STAGE_LUT[648] = -16'd104;
assign W_I_STAGE_LUT[648] = -16'd234;
assign W_R_STAGE_LUT[649] = -16'd104;
assign W_I_STAGE_LUT[649] = -16'd234;
assign W_R_STAGE_LUT[650] = -16'd105;
assign W_I_STAGE_LUT[650] = -16'd233;
assign W_R_STAGE_LUT[651] = -16'd106;
assign W_I_STAGE_LUT[651] = -16'd233;
assign W_R_STAGE_LUT[652] = -16'd107;
assign W_I_STAGE_LUT[652] = -16'd233;
assign W_R_STAGE_LUT[653] = -16'd107;
assign W_I_STAGE_LUT[653] = -16'd232;
assign W_R_STAGE_LUT[654] = -16'd108;
assign W_I_STAGE_LUT[654] = -16'd232;
assign W_R_STAGE_LUT[655] = -16'd109;
assign W_I_STAGE_LUT[655] = -16'd232;
assign W_R_STAGE_LUT[656] = -16'd109;
assign W_I_STAGE_LUT[656] = -16'd231;
assign W_R_STAGE_LUT[657] = -16'd110;
assign W_I_STAGE_LUT[657] = -16'd231;
assign W_R_STAGE_LUT[658] = -16'd111;
assign W_I_STAGE_LUT[658] = -16'd231;
assign W_R_STAGE_LUT[659] = -16'd112;
assign W_I_STAGE_LUT[659] = -16'd230;
assign W_R_STAGE_LUT[660] = -16'd112;
assign W_I_STAGE_LUT[660] = -16'd230;
assign W_R_STAGE_LUT[661] = -16'd113;
assign W_I_STAGE_LUT[661] = -16'd230;
assign W_R_STAGE_LUT[662] = -16'd114;
assign W_I_STAGE_LUT[662] = -16'd229;
assign W_R_STAGE_LUT[663] = -16'd114;
assign W_I_STAGE_LUT[663] = -16'd229;
assign W_R_STAGE_LUT[664] = -16'd115;
assign W_I_STAGE_LUT[664] = -16'd229;
assign W_R_STAGE_LUT[665] = -16'd116;
assign W_I_STAGE_LUT[665] = -16'd228;
assign W_R_STAGE_LUT[666] = -16'd117;
assign W_I_STAGE_LUT[666] = -16'd228;
assign W_R_STAGE_LUT[667] = -16'd117;
assign W_I_STAGE_LUT[667] = -16'd228;
assign W_R_STAGE_LUT[668] = -16'd118;
assign W_I_STAGE_LUT[668] = -16'd227;
assign W_R_STAGE_LUT[669] = -16'd119;
assign W_I_STAGE_LUT[669] = -16'd227;
assign W_R_STAGE_LUT[670] = -16'd119;
assign W_I_STAGE_LUT[670] = -16'd227;
assign W_R_STAGE_LUT[671] = -16'd120;
assign W_I_STAGE_LUT[671] = -16'd226;
assign W_R_STAGE_LUT[672] = -16'd121;
assign W_I_STAGE_LUT[672] = -16'd226;
assign W_R_STAGE_LUT[673] = -16'd121;
assign W_I_STAGE_LUT[673] = -16'd225;
assign W_R_STAGE_LUT[674] = -16'd122;
assign W_I_STAGE_LUT[674] = -16'd225;
assign W_R_STAGE_LUT[675] = -16'd123;
assign W_I_STAGE_LUT[675] = -16'd225;
assign W_R_STAGE_LUT[676] = -16'd123;
assign W_I_STAGE_LUT[676] = -16'd224;
assign W_R_STAGE_LUT[677] = -16'd124;
assign W_I_STAGE_LUT[677] = -16'd224;
assign W_R_STAGE_LUT[678] = -16'd125;
assign W_I_STAGE_LUT[678] = -16'd224;
assign W_R_STAGE_LUT[679] = -16'd125;
assign W_I_STAGE_LUT[679] = -16'd223;
assign W_R_STAGE_LUT[680] = -16'd126;
assign W_I_STAGE_LUT[680] = -16'd223;
assign W_R_STAGE_LUT[681] = -16'd127;
assign W_I_STAGE_LUT[681] = -16'd222;
assign W_R_STAGE_LUT[682] = -16'd128;
assign W_I_STAGE_LUT[682] = -16'd222;
assign W_R_STAGE_LUT[683] = -16'd128;
assign W_I_STAGE_LUT[683] = -16'd222;
assign W_R_STAGE_LUT[684] = -16'd129;
assign W_I_STAGE_LUT[684] = -16'd221;
assign W_R_STAGE_LUT[685] = -16'd130;
assign W_I_STAGE_LUT[685] = -16'd221;
assign W_R_STAGE_LUT[686] = -16'd130;
assign W_I_STAGE_LUT[686] = -16'd220;
assign W_R_STAGE_LUT[687] = -16'd131;
assign W_I_STAGE_LUT[687] = -16'd220;
assign W_R_STAGE_LUT[688] = -16'd132;
assign W_I_STAGE_LUT[688] = -16'd220;
assign W_R_STAGE_LUT[689] = -16'd132;
assign W_I_STAGE_LUT[689] = -16'd219;
assign W_R_STAGE_LUT[690] = -16'd133;
assign W_I_STAGE_LUT[690] = -16'd219;
assign W_R_STAGE_LUT[691] = -16'd134;
assign W_I_STAGE_LUT[691] = -16'd218;
assign W_R_STAGE_LUT[692] = -16'd134;
assign W_I_STAGE_LUT[692] = -16'd218;
assign W_R_STAGE_LUT[693] = -16'd135;
assign W_I_STAGE_LUT[693] = -16'd218;
assign W_R_STAGE_LUT[694] = -16'd136;
assign W_I_STAGE_LUT[694] = -16'd217;
assign W_R_STAGE_LUT[695] = -16'd136;
assign W_I_STAGE_LUT[695] = -16'd217;
assign W_R_STAGE_LUT[696] = -16'd137;
assign W_I_STAGE_LUT[696] = -16'd216;
assign W_R_STAGE_LUT[697] = -16'd138;
assign W_I_STAGE_LUT[697] = -16'd216;
assign W_R_STAGE_LUT[698] = -16'd138;
assign W_I_STAGE_LUT[698] = -16'd215;
assign W_R_STAGE_LUT[699] = -16'd139;
assign W_I_STAGE_LUT[699] = -16'd215;
assign W_R_STAGE_LUT[700] = -16'd140;
assign W_I_STAGE_LUT[700] = -16'd215;
assign W_R_STAGE_LUT[701] = -16'd140;
assign W_I_STAGE_LUT[701] = -16'd214;
assign W_R_STAGE_LUT[702] = -16'd141;
assign W_I_STAGE_LUT[702] = -16'd214;
assign W_R_STAGE_LUT[703] = -16'd142;
assign W_I_STAGE_LUT[703] = -16'd213;
assign W_R_STAGE_LUT[704] = -16'd142;
assign W_I_STAGE_LUT[704] = -16'd213;
assign W_R_STAGE_LUT[705] = -16'd143;
assign W_I_STAGE_LUT[705] = -16'd212;
assign W_R_STAGE_LUT[706] = -16'd144;
assign W_I_STAGE_LUT[706] = -16'd212;
assign W_R_STAGE_LUT[707] = -16'd144;
assign W_I_STAGE_LUT[707] = -16'd212;
assign W_R_STAGE_LUT[708] = -16'd145;
assign W_I_STAGE_LUT[708] = -16'd211;
assign W_R_STAGE_LUT[709] = -16'd145;
assign W_I_STAGE_LUT[709] = -16'd211;
assign W_R_STAGE_LUT[710] = -16'd146;
assign W_I_STAGE_LUT[710] = -16'd210;
assign W_R_STAGE_LUT[711] = -16'd147;
assign W_I_STAGE_LUT[711] = -16'd210;
assign W_R_STAGE_LUT[712] = -16'd147;
assign W_I_STAGE_LUT[712] = -16'd209;
assign W_R_STAGE_LUT[713] = -16'd148;
assign W_I_STAGE_LUT[713] = -16'd209;
assign W_R_STAGE_LUT[714] = -16'd149;
assign W_I_STAGE_LUT[714] = -16'd208;
assign W_R_STAGE_LUT[715] = -16'd149;
assign W_I_STAGE_LUT[715] = -16'd208;
assign W_R_STAGE_LUT[716] = -16'd150;
assign W_I_STAGE_LUT[716] = -16'd207;
assign W_R_STAGE_LUT[717] = -16'd151;
assign W_I_STAGE_LUT[717] = -16'd207;
assign W_R_STAGE_LUT[718] = -16'd151;
assign W_I_STAGE_LUT[718] = -16'd207;
assign W_R_STAGE_LUT[719] = -16'd152;
assign W_I_STAGE_LUT[719] = -16'd206;
assign W_R_STAGE_LUT[720] = -16'd152;
assign W_I_STAGE_LUT[720] = -16'd206;
assign W_R_STAGE_LUT[721] = -16'd153;
assign W_I_STAGE_LUT[721] = -16'd205;
assign W_R_STAGE_LUT[722] = -16'd154;
assign W_I_STAGE_LUT[722] = -16'd205;
assign W_R_STAGE_LUT[723] = -16'd154;
assign W_I_STAGE_LUT[723] = -16'd204;
assign W_R_STAGE_LUT[724] = -16'd155;
assign W_I_STAGE_LUT[724] = -16'd204;
assign W_R_STAGE_LUT[725] = -16'd156;
assign W_I_STAGE_LUT[725] = -16'd203;
assign W_R_STAGE_LUT[726] = -16'd156;
assign W_I_STAGE_LUT[726] = -16'd203;
assign W_R_STAGE_LUT[727] = -16'd157;
assign W_I_STAGE_LUT[727] = -16'd202;
assign W_R_STAGE_LUT[728] = -16'd157;
assign W_I_STAGE_LUT[728] = -16'd202;
assign W_R_STAGE_LUT[729] = -16'd158;
assign W_I_STAGE_LUT[729] = -16'd201;
assign W_R_STAGE_LUT[730] = -16'd159;
assign W_I_STAGE_LUT[730] = -16'd201;
assign W_R_STAGE_LUT[731] = -16'd159;
assign W_I_STAGE_LUT[731] = -16'd200;
assign W_R_STAGE_LUT[732] = -16'd160;
assign W_I_STAGE_LUT[732] = -16'd200;
assign W_R_STAGE_LUT[733] = -16'd161;
assign W_I_STAGE_LUT[733] = -16'd199;
assign W_R_STAGE_LUT[734] = -16'd161;
assign W_I_STAGE_LUT[734] = -16'd199;
assign W_R_STAGE_LUT[735] = -16'd162;
assign W_I_STAGE_LUT[735] = -16'd198;
assign W_R_STAGE_LUT[736] = -16'd162;
assign W_I_STAGE_LUT[736] = -16'd198;
assign W_R_STAGE_LUT[737] = -16'd163;
assign W_I_STAGE_LUT[737] = -16'd197;
assign W_R_STAGE_LUT[738] = -16'd164;
assign W_I_STAGE_LUT[738] = -16'd197;
assign W_R_STAGE_LUT[739] = -16'd164;
assign W_I_STAGE_LUT[739] = -16'd196;
assign W_R_STAGE_LUT[740] = -16'd165;
assign W_I_STAGE_LUT[740] = -16'd196;
assign W_R_STAGE_LUT[741] = -16'd165;
assign W_I_STAGE_LUT[741] = -16'd195;
assign W_R_STAGE_LUT[742] = -16'd166;
assign W_I_STAGE_LUT[742] = -16'd195;
assign W_R_STAGE_LUT[743] = -16'd167;
assign W_I_STAGE_LUT[743] = -16'd194;
assign W_R_STAGE_LUT[744] = -16'd167;
assign W_I_STAGE_LUT[744] = -16'd194;
assign W_R_STAGE_LUT[745] = -16'd168;
assign W_I_STAGE_LUT[745] = -16'd193;
assign W_R_STAGE_LUT[746] = -16'd168;
assign W_I_STAGE_LUT[746] = -16'd193;
assign W_R_STAGE_LUT[747] = -16'd169;
assign W_I_STAGE_LUT[747] = -16'd192;
assign W_R_STAGE_LUT[748] = -16'd170;
assign W_I_STAGE_LUT[748] = -16'd192;
assign W_R_STAGE_LUT[749] = -16'd170;
assign W_I_STAGE_LUT[749] = -16'd191;
assign W_R_STAGE_LUT[750] = -16'd171;
assign W_I_STAGE_LUT[750] = -16'd191;
assign W_R_STAGE_LUT[751] = -16'd171;
assign W_I_STAGE_LUT[751] = -16'd190;
assign W_R_STAGE_LUT[752] = -16'd172;
assign W_I_STAGE_LUT[752] = -16'd190;
assign W_R_STAGE_LUT[753] = -16'd173;
assign W_I_STAGE_LUT[753] = -16'd189;
assign W_R_STAGE_LUT[754] = -16'd173;
assign W_I_STAGE_LUT[754] = -16'd189;
assign W_R_STAGE_LUT[755] = -16'd174;
assign W_I_STAGE_LUT[755] = -16'd188;
assign W_R_STAGE_LUT[756] = -16'd174;
assign W_I_STAGE_LUT[756] = -16'd188;
assign W_R_STAGE_LUT[757] = -16'd175;
assign W_I_STAGE_LUT[757] = -16'd187;
assign W_R_STAGE_LUT[758] = -16'd175;
assign W_I_STAGE_LUT[758] = -16'd186;
assign W_R_STAGE_LUT[759] = -16'd176;
assign W_I_STAGE_LUT[759] = -16'd186;
assign W_R_STAGE_LUT[760] = -16'd177;
assign W_I_STAGE_LUT[760] = -16'd185;
assign W_R_STAGE_LUT[761] = -16'd177;
assign W_I_STAGE_LUT[761] = -16'd185;
assign W_R_STAGE_LUT[762] = -16'd178;
assign W_I_STAGE_LUT[762] = -16'd184;
assign W_R_STAGE_LUT[763] = -16'd178;
assign W_I_STAGE_LUT[763] = -16'd184;
assign W_R_STAGE_LUT[764] = -16'd179;
assign W_I_STAGE_LUT[764] = -16'd183;
assign W_R_STAGE_LUT[765] = -16'd179;
assign W_I_STAGE_LUT[765] = -16'd183;
assign W_R_STAGE_LUT[766] = -16'd180;
assign W_I_STAGE_LUT[766] = -16'd182;
assign W_R_STAGE_LUT[767] = -16'd180;
assign W_I_STAGE_LUT[767] = -16'd182;
assign W_R_STAGE_LUT[768] = -16'd181;
assign W_I_STAGE_LUT[768] = -16'd181;
assign W_R_STAGE_LUT[769] = -16'd182;
assign W_I_STAGE_LUT[769] = -16'd180;
assign W_R_STAGE_LUT[770] = -16'd182;
assign W_I_STAGE_LUT[770] = -16'd180;
assign W_R_STAGE_LUT[771] = -16'd183;
assign W_I_STAGE_LUT[771] = -16'd179;
assign W_R_STAGE_LUT[772] = -16'd183;
assign W_I_STAGE_LUT[772] = -16'd179;
assign W_R_STAGE_LUT[773] = -16'd184;
assign W_I_STAGE_LUT[773] = -16'd178;
assign W_R_STAGE_LUT[774] = -16'd184;
assign W_I_STAGE_LUT[774] = -16'd178;
assign W_R_STAGE_LUT[775] = -16'd185;
assign W_I_STAGE_LUT[775] = -16'd177;
assign W_R_STAGE_LUT[776] = -16'd185;
assign W_I_STAGE_LUT[776] = -16'd177;
assign W_R_STAGE_LUT[777] = -16'd186;
assign W_I_STAGE_LUT[777] = -16'd176;
assign W_R_STAGE_LUT[778] = -16'd186;
assign W_I_STAGE_LUT[778] = -16'd175;
assign W_R_STAGE_LUT[779] = -16'd187;
assign W_I_STAGE_LUT[779] = -16'd175;
assign W_R_STAGE_LUT[780] = -16'd188;
assign W_I_STAGE_LUT[780] = -16'd174;
assign W_R_STAGE_LUT[781] = -16'd188;
assign W_I_STAGE_LUT[781] = -16'd174;
assign W_R_STAGE_LUT[782] = -16'd189;
assign W_I_STAGE_LUT[782] = -16'd173;
assign W_R_STAGE_LUT[783] = -16'd189;
assign W_I_STAGE_LUT[783] = -16'd173;
assign W_R_STAGE_LUT[784] = -16'd190;
assign W_I_STAGE_LUT[784] = -16'd172;
assign W_R_STAGE_LUT[785] = -16'd190;
assign W_I_STAGE_LUT[785] = -16'd171;
assign W_R_STAGE_LUT[786] = -16'd191;
assign W_I_STAGE_LUT[786] = -16'd171;
assign W_R_STAGE_LUT[787] = -16'd191;
assign W_I_STAGE_LUT[787] = -16'd170;
assign W_R_STAGE_LUT[788] = -16'd192;
assign W_I_STAGE_LUT[788] = -16'd170;
assign W_R_STAGE_LUT[789] = -16'd192;
assign W_I_STAGE_LUT[789] = -16'd169;
assign W_R_STAGE_LUT[790] = -16'd193;
assign W_I_STAGE_LUT[790] = -16'd168;
assign W_R_STAGE_LUT[791] = -16'd193;
assign W_I_STAGE_LUT[791] = -16'd168;
assign W_R_STAGE_LUT[792] = -16'd194;
assign W_I_STAGE_LUT[792] = -16'd167;
assign W_R_STAGE_LUT[793] = -16'd194;
assign W_I_STAGE_LUT[793] = -16'd167;
assign W_R_STAGE_LUT[794] = -16'd195;
assign W_I_STAGE_LUT[794] = -16'd166;
assign W_R_STAGE_LUT[795] = -16'd195;
assign W_I_STAGE_LUT[795] = -16'd165;
assign W_R_STAGE_LUT[796] = -16'd196;
assign W_I_STAGE_LUT[796] = -16'd165;
assign W_R_STAGE_LUT[797] = -16'd196;
assign W_I_STAGE_LUT[797] = -16'd164;
assign W_R_STAGE_LUT[798] = -16'd197;
assign W_I_STAGE_LUT[798] = -16'd164;
assign W_R_STAGE_LUT[799] = -16'd197;
assign W_I_STAGE_LUT[799] = -16'd163;
assign W_R_STAGE_LUT[800] = -16'd198;
assign W_I_STAGE_LUT[800] = -16'd162;
assign W_R_STAGE_LUT[801] = -16'd198;
assign W_I_STAGE_LUT[801] = -16'd162;
assign W_R_STAGE_LUT[802] = -16'd199;
assign W_I_STAGE_LUT[802] = -16'd161;
assign W_R_STAGE_LUT[803] = -16'd199;
assign W_I_STAGE_LUT[803] = -16'd161;
assign W_R_STAGE_LUT[804] = -16'd200;
assign W_I_STAGE_LUT[804] = -16'd160;
assign W_R_STAGE_LUT[805] = -16'd200;
assign W_I_STAGE_LUT[805] = -16'd159;
assign W_R_STAGE_LUT[806] = -16'd201;
assign W_I_STAGE_LUT[806] = -16'd159;
assign W_R_STAGE_LUT[807] = -16'd201;
assign W_I_STAGE_LUT[807] = -16'd158;
assign W_R_STAGE_LUT[808] = -16'd202;
assign W_I_STAGE_LUT[808] = -16'd157;
assign W_R_STAGE_LUT[809] = -16'd202;
assign W_I_STAGE_LUT[809] = -16'd157;
assign W_R_STAGE_LUT[810] = -16'd203;
assign W_I_STAGE_LUT[810] = -16'd156;
assign W_R_STAGE_LUT[811] = -16'd203;
assign W_I_STAGE_LUT[811] = -16'd156;
assign W_R_STAGE_LUT[812] = -16'd204;
assign W_I_STAGE_LUT[812] = -16'd155;
assign W_R_STAGE_LUT[813] = -16'd204;
assign W_I_STAGE_LUT[813] = -16'd154;
assign W_R_STAGE_LUT[814] = -16'd205;
assign W_I_STAGE_LUT[814] = -16'd154;
assign W_R_STAGE_LUT[815] = -16'd205;
assign W_I_STAGE_LUT[815] = -16'd153;
assign W_R_STAGE_LUT[816] = -16'd206;
assign W_I_STAGE_LUT[816] = -16'd152;
assign W_R_STAGE_LUT[817] = -16'd206;
assign W_I_STAGE_LUT[817] = -16'd152;
assign W_R_STAGE_LUT[818] = -16'd207;
assign W_I_STAGE_LUT[818] = -16'd151;
assign W_R_STAGE_LUT[819] = -16'd207;
assign W_I_STAGE_LUT[819] = -16'd151;
assign W_R_STAGE_LUT[820] = -16'd207;
assign W_I_STAGE_LUT[820] = -16'd150;
assign W_R_STAGE_LUT[821] = -16'd208;
assign W_I_STAGE_LUT[821] = -16'd149;
assign W_R_STAGE_LUT[822] = -16'd208;
assign W_I_STAGE_LUT[822] = -16'd149;
assign W_R_STAGE_LUT[823] = -16'd209;
assign W_I_STAGE_LUT[823] = -16'd148;
assign W_R_STAGE_LUT[824] = -16'd209;
assign W_I_STAGE_LUT[824] = -16'd147;
assign W_R_STAGE_LUT[825] = -16'd210;
assign W_I_STAGE_LUT[825] = -16'd147;
assign W_R_STAGE_LUT[826] = -16'd210;
assign W_I_STAGE_LUT[826] = -16'd146;
assign W_R_STAGE_LUT[827] = -16'd211;
assign W_I_STAGE_LUT[827] = -16'd145;
assign W_R_STAGE_LUT[828] = -16'd211;
assign W_I_STAGE_LUT[828] = -16'd145;
assign W_R_STAGE_LUT[829] = -16'd212;
assign W_I_STAGE_LUT[829] = -16'd144;
assign W_R_STAGE_LUT[830] = -16'd212;
assign W_I_STAGE_LUT[830] = -16'd144;
assign W_R_STAGE_LUT[831] = -16'd212;
assign W_I_STAGE_LUT[831] = -16'd143;
assign W_R_STAGE_LUT[832] = -16'd213;
assign W_I_STAGE_LUT[832] = -16'd142;
assign W_R_STAGE_LUT[833] = -16'd213;
assign W_I_STAGE_LUT[833] = -16'd142;
assign W_R_STAGE_LUT[834] = -16'd214;
assign W_I_STAGE_LUT[834] = -16'd141;
assign W_R_STAGE_LUT[835] = -16'd214;
assign W_I_STAGE_LUT[835] = -16'd140;
assign W_R_STAGE_LUT[836] = -16'd215;
assign W_I_STAGE_LUT[836] = -16'd140;
assign W_R_STAGE_LUT[837] = -16'd215;
assign W_I_STAGE_LUT[837] = -16'd139;
assign W_R_STAGE_LUT[838] = -16'd215;
assign W_I_STAGE_LUT[838] = -16'd138;
assign W_R_STAGE_LUT[839] = -16'd216;
assign W_I_STAGE_LUT[839] = -16'd138;
assign W_R_STAGE_LUT[840] = -16'd216;
assign W_I_STAGE_LUT[840] = -16'd137;
assign W_R_STAGE_LUT[841] = -16'd217;
assign W_I_STAGE_LUT[841] = -16'd136;
assign W_R_STAGE_LUT[842] = -16'd217;
assign W_I_STAGE_LUT[842] = -16'd136;
assign W_R_STAGE_LUT[843] = -16'd218;
assign W_I_STAGE_LUT[843] = -16'd135;
assign W_R_STAGE_LUT[844] = -16'd218;
assign W_I_STAGE_LUT[844] = -16'd134;
assign W_R_STAGE_LUT[845] = -16'd218;
assign W_I_STAGE_LUT[845] = -16'd134;
assign W_R_STAGE_LUT[846] = -16'd219;
assign W_I_STAGE_LUT[846] = -16'd133;
assign W_R_STAGE_LUT[847] = -16'd219;
assign W_I_STAGE_LUT[847] = -16'd132;
assign W_R_STAGE_LUT[848] = -16'd220;
assign W_I_STAGE_LUT[848] = -16'd132;
assign W_R_STAGE_LUT[849] = -16'd220;
assign W_I_STAGE_LUT[849] = -16'd131;
assign W_R_STAGE_LUT[850] = -16'd220;
assign W_I_STAGE_LUT[850] = -16'd130;
assign W_R_STAGE_LUT[851] = -16'd221;
assign W_I_STAGE_LUT[851] = -16'd130;
assign W_R_STAGE_LUT[852] = -16'd221;
assign W_I_STAGE_LUT[852] = -16'd129;
assign W_R_STAGE_LUT[853] = -16'd222;
assign W_I_STAGE_LUT[853] = -16'd128;
assign W_R_STAGE_LUT[854] = -16'd222;
assign W_I_STAGE_LUT[854] = -16'd128;
assign W_R_STAGE_LUT[855] = -16'd222;
assign W_I_STAGE_LUT[855] = -16'd127;
assign W_R_STAGE_LUT[856] = -16'd223;
assign W_I_STAGE_LUT[856] = -16'd126;
assign W_R_STAGE_LUT[857] = -16'd223;
assign W_I_STAGE_LUT[857] = -16'd125;
assign W_R_STAGE_LUT[858] = -16'd224;
assign W_I_STAGE_LUT[858] = -16'd125;
assign W_R_STAGE_LUT[859] = -16'd224;
assign W_I_STAGE_LUT[859] = -16'd124;
assign W_R_STAGE_LUT[860] = -16'd224;
assign W_I_STAGE_LUT[860] = -16'd123;
assign W_R_STAGE_LUT[861] = -16'd225;
assign W_I_STAGE_LUT[861] = -16'd123;
assign W_R_STAGE_LUT[862] = -16'd225;
assign W_I_STAGE_LUT[862] = -16'd122;
assign W_R_STAGE_LUT[863] = -16'd225;
assign W_I_STAGE_LUT[863] = -16'd121;
assign W_R_STAGE_LUT[864] = -16'd226;
assign W_I_STAGE_LUT[864] = -16'd121;
assign W_R_STAGE_LUT[865] = -16'd226;
assign W_I_STAGE_LUT[865] = -16'd120;
assign W_R_STAGE_LUT[866] = -16'd227;
assign W_I_STAGE_LUT[866] = -16'd119;
assign W_R_STAGE_LUT[867] = -16'd227;
assign W_I_STAGE_LUT[867] = -16'd119;
assign W_R_STAGE_LUT[868] = -16'd227;
assign W_I_STAGE_LUT[868] = -16'd118;
assign W_R_STAGE_LUT[869] = -16'd228;
assign W_I_STAGE_LUT[869] = -16'd117;
assign W_R_STAGE_LUT[870] = -16'd228;
assign W_I_STAGE_LUT[870] = -16'd117;
assign W_R_STAGE_LUT[871] = -16'd228;
assign W_I_STAGE_LUT[871] = -16'd116;
assign W_R_STAGE_LUT[872] = -16'd229;
assign W_I_STAGE_LUT[872] = -16'd115;
assign W_R_STAGE_LUT[873] = -16'd229;
assign W_I_STAGE_LUT[873] = -16'd114;
assign W_R_STAGE_LUT[874] = -16'd229;
assign W_I_STAGE_LUT[874] = -16'd114;
assign W_R_STAGE_LUT[875] = -16'd230;
assign W_I_STAGE_LUT[875] = -16'd113;
assign W_R_STAGE_LUT[876] = -16'd230;
assign W_I_STAGE_LUT[876] = -16'd112;
assign W_R_STAGE_LUT[877] = -16'd230;
assign W_I_STAGE_LUT[877] = -16'd112;
assign W_R_STAGE_LUT[878] = -16'd231;
assign W_I_STAGE_LUT[878] = -16'd111;
assign W_R_STAGE_LUT[879] = -16'd231;
assign W_I_STAGE_LUT[879] = -16'd110;
assign W_R_STAGE_LUT[880] = -16'd231;
assign W_I_STAGE_LUT[880] = -16'd109;
assign W_R_STAGE_LUT[881] = -16'd232;
assign W_I_STAGE_LUT[881] = -16'd109;
assign W_R_STAGE_LUT[882] = -16'd232;
assign W_I_STAGE_LUT[882] = -16'd108;
assign W_R_STAGE_LUT[883] = -16'd232;
assign W_I_STAGE_LUT[883] = -16'd107;
assign W_R_STAGE_LUT[884] = -16'd233;
assign W_I_STAGE_LUT[884] = -16'd107;
assign W_R_STAGE_LUT[885] = -16'd233;
assign W_I_STAGE_LUT[885] = -16'd106;
assign W_R_STAGE_LUT[886] = -16'd233;
assign W_I_STAGE_LUT[886] = -16'd105;
assign W_R_STAGE_LUT[887] = -16'd234;
assign W_I_STAGE_LUT[887] = -16'd104;
assign W_R_STAGE_LUT[888] = -16'd234;
assign W_I_STAGE_LUT[888] = -16'd104;
assign W_R_STAGE_LUT[889] = -16'd234;
assign W_I_STAGE_LUT[889] = -16'd103;
assign W_R_STAGE_LUT[890] = -16'd235;
assign W_I_STAGE_LUT[890] = -16'd102;
assign W_R_STAGE_LUT[891] = -16'd235;
assign W_I_STAGE_LUT[891] = -16'd102;
assign W_R_STAGE_LUT[892] = -16'd235;
assign W_I_STAGE_LUT[892] = -16'd101;
assign W_R_STAGE_LUT[893] = -16'd236;
assign W_I_STAGE_LUT[893] = -16'd100;
assign W_R_STAGE_LUT[894] = -16'd236;
assign W_I_STAGE_LUT[894] = -16'd99;
assign W_R_STAGE_LUT[895] = -16'd236;
assign W_I_STAGE_LUT[895] = -16'd99;
assign W_R_STAGE_LUT[896] = -16'd237;
assign W_I_STAGE_LUT[896] = -16'd98;
assign W_R_STAGE_LUT[897] = -16'd237;
assign W_I_STAGE_LUT[897] = -16'd97;
assign W_R_STAGE_LUT[898] = -16'd237;
assign W_I_STAGE_LUT[898] = -16'd97;
assign W_R_STAGE_LUT[899] = -16'd237;
assign W_I_STAGE_LUT[899] = -16'd96;
assign W_R_STAGE_LUT[900] = -16'd238;
assign W_I_STAGE_LUT[900] = -16'd95;
assign W_R_STAGE_LUT[901] = -16'd238;
assign W_I_STAGE_LUT[901] = -16'd94;
assign W_R_STAGE_LUT[902] = -16'd238;
assign W_I_STAGE_LUT[902] = -16'd94;
assign W_R_STAGE_LUT[903] = -16'd239;
assign W_I_STAGE_LUT[903] = -16'd93;
assign W_R_STAGE_LUT[904] = -16'd239;
assign W_I_STAGE_LUT[904] = -16'd92;
assign W_R_STAGE_LUT[905] = -16'd239;
assign W_I_STAGE_LUT[905] = -16'd91;
assign W_R_STAGE_LUT[906] = -16'd239;
assign W_I_STAGE_LUT[906] = -16'd91;
assign W_R_STAGE_LUT[907] = -16'd240;
assign W_I_STAGE_LUT[907] = -16'd90;
assign W_R_STAGE_LUT[908] = -16'd240;
assign W_I_STAGE_LUT[908] = -16'd89;
assign W_R_STAGE_LUT[909] = -16'd240;
assign W_I_STAGE_LUT[909] = -16'd88;
assign W_R_STAGE_LUT[910] = -16'd241;
assign W_I_STAGE_LUT[910] = -16'd88;
assign W_R_STAGE_LUT[911] = -16'd241;
assign W_I_STAGE_LUT[911] = -16'd87;
assign W_R_STAGE_LUT[912] = -16'd241;
assign W_I_STAGE_LUT[912] = -16'd86;
assign W_R_STAGE_LUT[913] = -16'd241;
assign W_I_STAGE_LUT[913] = -16'd86;
assign W_R_STAGE_LUT[914] = -16'd242;
assign W_I_STAGE_LUT[914] = -16'd85;
assign W_R_STAGE_LUT[915] = -16'd242;
assign W_I_STAGE_LUT[915] = -16'd84;
assign W_R_STAGE_LUT[916] = -16'd242;
assign W_I_STAGE_LUT[916] = -16'd83;
assign W_R_STAGE_LUT[917] = -16'd242;
assign W_I_STAGE_LUT[917] = -16'd83;
assign W_R_STAGE_LUT[918] = -16'd243;
assign W_I_STAGE_LUT[918] = -16'd82;
assign W_R_STAGE_LUT[919] = -16'd243;
assign W_I_STAGE_LUT[919] = -16'd81;
assign W_R_STAGE_LUT[920] = -16'd243;
assign W_I_STAGE_LUT[920] = -16'd80;
assign W_R_STAGE_LUT[921] = -16'd243;
assign W_I_STAGE_LUT[921] = -16'd80;
assign W_R_STAGE_LUT[922] = -16'd244;
assign W_I_STAGE_LUT[922] = -16'd79;
assign W_R_STAGE_LUT[923] = -16'd244;
assign W_I_STAGE_LUT[923] = -16'd78;
assign W_R_STAGE_LUT[924] = -16'd244;
assign W_I_STAGE_LUT[924] = -16'd77;
assign W_R_STAGE_LUT[925] = -16'd244;
assign W_I_STAGE_LUT[925] = -16'd77;
assign W_R_STAGE_LUT[926] = -16'd245;
assign W_I_STAGE_LUT[926] = -16'd76;
assign W_R_STAGE_LUT[927] = -16'd245;
assign W_I_STAGE_LUT[927] = -16'd75;
assign W_R_STAGE_LUT[928] = -16'd245;
assign W_I_STAGE_LUT[928] = -16'd74;
assign W_R_STAGE_LUT[929] = -16'd245;
assign W_I_STAGE_LUT[929] = -16'd74;
assign W_R_STAGE_LUT[930] = -16'd245;
assign W_I_STAGE_LUT[930] = -16'd73;
assign W_R_STAGE_LUT[931] = -16'd246;
assign W_I_STAGE_LUT[931] = -16'd72;
assign W_R_STAGE_LUT[932] = -16'd246;
assign W_I_STAGE_LUT[932] = -16'd71;
assign W_R_STAGE_LUT[933] = -16'd246;
assign W_I_STAGE_LUT[933] = -16'd71;
assign W_R_STAGE_LUT[934] = -16'd246;
assign W_I_STAGE_LUT[934] = -16'd70;
assign W_R_STAGE_LUT[935] = -16'd247;
assign W_I_STAGE_LUT[935] = -16'd69;
assign W_R_STAGE_LUT[936] = -16'd247;
assign W_I_STAGE_LUT[936] = -16'd68;
assign W_R_STAGE_LUT[937] = -16'd247;
assign W_I_STAGE_LUT[937] = -16'd68;
assign W_R_STAGE_LUT[938] = -16'd247;
assign W_I_STAGE_LUT[938] = -16'd67;
assign W_R_STAGE_LUT[939] = -16'd247;
assign W_I_STAGE_LUT[939] = -16'd66;
assign W_R_STAGE_LUT[940] = -16'd248;
assign W_I_STAGE_LUT[940] = -16'd65;
assign W_R_STAGE_LUT[941] = -16'd248;
assign W_I_STAGE_LUT[941] = -16'd64;
assign W_R_STAGE_LUT[942] = -16'd248;
assign W_I_STAGE_LUT[942] = -16'd64;
assign W_R_STAGE_LUT[943] = -16'd248;
assign W_I_STAGE_LUT[943] = -16'd63;
assign W_R_STAGE_LUT[944] = -16'd248;
assign W_I_STAGE_LUT[944] = -16'd62;
assign W_R_STAGE_LUT[945] = -16'd249;
assign W_I_STAGE_LUT[945] = -16'd61;
assign W_R_STAGE_LUT[946] = -16'd249;
assign W_I_STAGE_LUT[946] = -16'd61;
assign W_R_STAGE_LUT[947] = -16'd249;
assign W_I_STAGE_LUT[947] = -16'd60;
assign W_R_STAGE_LUT[948] = -16'd249;
assign W_I_STAGE_LUT[948] = -16'd59;
assign W_R_STAGE_LUT[949] = -16'd249;
assign W_I_STAGE_LUT[949] = -16'd58;
assign W_R_STAGE_LUT[950] = -16'd249;
assign W_I_STAGE_LUT[950] = -16'd58;
assign W_R_STAGE_LUT[951] = -16'd250;
assign W_I_STAGE_LUT[951] = -16'd57;
assign W_R_STAGE_LUT[952] = -16'd250;
assign W_I_STAGE_LUT[952] = -16'd56;
assign W_R_STAGE_LUT[953] = -16'd250;
assign W_I_STAGE_LUT[953] = -16'd55;
assign W_R_STAGE_LUT[954] = -16'd250;
assign W_I_STAGE_LUT[954] = -16'd55;
assign W_R_STAGE_LUT[955] = -16'd250;
assign W_I_STAGE_LUT[955] = -16'd54;
assign W_R_STAGE_LUT[956] = -16'd250;
assign W_I_STAGE_LUT[956] = -16'd53;
assign W_R_STAGE_LUT[957] = -16'd251;
assign W_I_STAGE_LUT[957] = -16'd52;
assign W_R_STAGE_LUT[958] = -16'd251;
assign W_I_STAGE_LUT[958] = -16'd51;
assign W_R_STAGE_LUT[959] = -16'd251;
assign W_I_STAGE_LUT[959] = -16'd51;
assign W_R_STAGE_LUT[960] = -16'd251;
assign W_I_STAGE_LUT[960] = -16'd50;
assign W_R_STAGE_LUT[961] = -16'd251;
assign W_I_STAGE_LUT[961] = -16'd49;
assign W_R_STAGE_LUT[962] = -16'd251;
assign W_I_STAGE_LUT[962] = -16'd48;
assign W_R_STAGE_LUT[963] = -16'd252;
assign W_I_STAGE_LUT[963] = -16'd48;
assign W_R_STAGE_LUT[964] = -16'd252;
assign W_I_STAGE_LUT[964] = -16'd47;
assign W_R_STAGE_LUT[965] = -16'd252;
assign W_I_STAGE_LUT[965] = -16'd46;
assign W_R_STAGE_LUT[966] = -16'd252;
assign W_I_STAGE_LUT[966] = -16'd45;
assign W_R_STAGE_LUT[967] = -16'd252;
assign W_I_STAGE_LUT[967] = -16'd45;
assign W_R_STAGE_LUT[968] = -16'd252;
assign W_I_STAGE_LUT[968] = -16'd44;
assign W_R_STAGE_LUT[969] = -16'd252;
assign W_I_STAGE_LUT[969] = -16'd43;
assign W_R_STAGE_LUT[970] = -16'd252;
assign W_I_STAGE_LUT[970] = -16'd42;
assign W_R_STAGE_LUT[971] = -16'd253;
assign W_I_STAGE_LUT[971] = -16'd41;
assign W_R_STAGE_LUT[972] = -16'd253;
assign W_I_STAGE_LUT[972] = -16'd41;
assign W_R_STAGE_LUT[973] = -16'd253;
assign W_I_STAGE_LUT[973] = -16'd40;
assign W_R_STAGE_LUT[974] = -16'd253;
assign W_I_STAGE_LUT[974] = -16'd39;
assign W_R_STAGE_LUT[975] = -16'd253;
assign W_I_STAGE_LUT[975] = -16'd38;
assign W_R_STAGE_LUT[976] = -16'd253;
assign W_I_STAGE_LUT[976] = -16'd38;
assign W_R_STAGE_LUT[977] = -16'd253;
assign W_I_STAGE_LUT[977] = -16'd37;
assign W_R_STAGE_LUT[978] = -16'd253;
assign W_I_STAGE_LUT[978] = -16'd36;
assign W_R_STAGE_LUT[979] = -16'd254;
assign W_I_STAGE_LUT[979] = -16'd35;
assign W_R_STAGE_LUT[980] = -16'd254;
assign W_I_STAGE_LUT[980] = -16'd34;
assign W_R_STAGE_LUT[981] = -16'd254;
assign W_I_STAGE_LUT[981] = -16'd34;
assign W_R_STAGE_LUT[982] = -16'd254;
assign W_I_STAGE_LUT[982] = -16'd33;
assign W_R_STAGE_LUT[983] = -16'd254;
assign W_I_STAGE_LUT[983] = -16'd32;
assign W_R_STAGE_LUT[984] = -16'd254;
assign W_I_STAGE_LUT[984] = -16'd31;
assign W_R_STAGE_LUT[985] = -16'd254;
assign W_I_STAGE_LUT[985] = -16'd31;
assign W_R_STAGE_LUT[986] = -16'd254;
assign W_I_STAGE_LUT[986] = -16'd30;
assign W_R_STAGE_LUT[987] = -16'd254;
assign W_I_STAGE_LUT[987] = -16'd29;
assign W_R_STAGE_LUT[988] = -16'd254;
assign W_I_STAGE_LUT[988] = -16'd28;
assign W_R_STAGE_LUT[989] = -16'd255;
assign W_I_STAGE_LUT[989] = -16'd27;
assign W_R_STAGE_LUT[990] = -16'd255;
assign W_I_STAGE_LUT[990] = -16'd27;
assign W_R_STAGE_LUT[991] = -16'd255;
assign W_I_STAGE_LUT[991] = -16'd26;
assign W_R_STAGE_LUT[992] = -16'd255;
assign W_I_STAGE_LUT[992] = -16'd25;
assign W_R_STAGE_LUT[993] = -16'd255;
assign W_I_STAGE_LUT[993] = -16'd24;
assign W_R_STAGE_LUT[994] = -16'd255;
assign W_I_STAGE_LUT[994] = -16'd24;
assign W_R_STAGE_LUT[995] = -16'd255;
assign W_I_STAGE_LUT[995] = -16'd23;
assign W_R_STAGE_LUT[996] = -16'd255;
assign W_I_STAGE_LUT[996] = -16'd22;
assign W_R_STAGE_LUT[997] = -16'd255;
assign W_I_STAGE_LUT[997] = -16'd21;
assign W_R_STAGE_LUT[998] = -16'd255;
assign W_I_STAGE_LUT[998] = -16'd20;
assign W_R_STAGE_LUT[999] = -16'd255;
assign W_I_STAGE_LUT[999] = -16'd20;
assign W_R_STAGE_LUT[1000] = -16'd255;
assign W_I_STAGE_LUT[1000] = -16'd19;
assign W_R_STAGE_LUT[1001] = -16'd255;
assign W_I_STAGE_LUT[1001] = -16'd18;
assign W_R_STAGE_LUT[1002] = -16'd255;
assign W_I_STAGE_LUT[1002] = -16'd17;
assign W_R_STAGE_LUT[1003] = -16'd255;
assign W_I_STAGE_LUT[1003] = -16'd16;
assign W_R_STAGE_LUT[1004] = -16'd256;
assign W_I_STAGE_LUT[1004] = -16'd16;
assign W_R_STAGE_LUT[1005] = -16'd256;
assign W_I_STAGE_LUT[1005] = -16'd15;
assign W_R_STAGE_LUT[1006] = -16'd256;
assign W_I_STAGE_LUT[1006] = -16'd14;
assign W_R_STAGE_LUT[1007] = -16'd256;
assign W_I_STAGE_LUT[1007] = -16'd13;
assign W_R_STAGE_LUT[1008] = -16'd256;
assign W_I_STAGE_LUT[1008] = -16'd13;
assign W_R_STAGE_LUT[1009] = -16'd256;
assign W_I_STAGE_LUT[1009] = -16'd12;
assign W_R_STAGE_LUT[1010] = -16'd256;
assign W_I_STAGE_LUT[1010] = -16'd11;
assign W_R_STAGE_LUT[1011] = -16'd256;
assign W_I_STAGE_LUT[1011] = -16'd10;
assign W_R_STAGE_LUT[1012] = -16'd256;
assign W_I_STAGE_LUT[1012] = -16'd9;
assign W_R_STAGE_LUT[1013] = -16'd256;
assign W_I_STAGE_LUT[1013] = -16'd9;
assign W_R_STAGE_LUT[1014] = -16'd256;
assign W_I_STAGE_LUT[1014] = -16'd8;
assign W_R_STAGE_LUT[1015] = -16'd256;
assign W_I_STAGE_LUT[1015] = -16'd7;
assign W_R_STAGE_LUT[1016] = -16'd256;
assign W_I_STAGE_LUT[1016] = -16'd6;
assign W_R_STAGE_LUT[1017] = -16'd256;
assign W_I_STAGE_LUT[1017] = -16'd5;
assign W_R_STAGE_LUT[1018] = -16'd256;
assign W_I_STAGE_LUT[1018] = -16'd5;
assign W_R_STAGE_LUT[1019] = -16'd256;
assign W_I_STAGE_LUT[1019] = -16'd4;
assign W_R_STAGE_LUT[1020] = -16'd256;
assign W_I_STAGE_LUT[1020] = -16'd3;
assign W_R_STAGE_LUT[1021] = -16'd256;
assign W_I_STAGE_LUT[1021] = -16'd2;
assign W_R_STAGE_LUT[1022] = -16'd256;
assign W_I_STAGE_LUT[1022] = -16'd2;
assign W_R_STAGE_LUT[1023] = -16'd256;
assign W_I_STAGE_LUT[1023] = -16'd1;
